* NGSPICE file created from fsm_flat.ext - technology: ihp-sg13g2

.subckt fsm_flat Timer_en adc_en clk_gating_en power_on sc_en timer_done tx_start
+ uart_busy uart_done uart_en adc_done adc_start clk reset wake_up_sg VDD VSS
N0 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=2.28077n ps=0.01084 w=0.42u l=1u
N1 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=3.17827n ps=0.01242 w=1u l=1u
N2 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N4 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N5 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N6 VSS a_16048_15454# a_15697_15311# VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
N7 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N8 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N9 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N10 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N11 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N12 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N13 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N14 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N15 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N16 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N17 a_14697_16043# a_14340_16000# VDD VDD sg13g2_lv_pmos ad=63f pd=0.72u as=0.1563p ps=1.22u w=0.42u l=0.13u
N18 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N19 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N20 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N21 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N22 a_14054_16434# sg13g2_inv_1_1.Y VDD VDD sg13g2_lv_pmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
N23 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N24 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N25 a_11654_13722# a_12459_13844# a_11914_13945# VDD sg13g2_lv_pmos ad=0.1428p pd=1.52u as=79.8f ps=0.8u w=0.42u l=0.13u
N26 VSS sg13g2_a21oi_1_0.A1 a_14248_23556# VSS sg13g2_lv_nmos ad=0.14875p pd=1.16u as=0.187p ps=1.78u w=0.55u l=0.13u
N27 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N28 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N29 VDD sg13g2_inv_1_0.Y a_12394_14452# VDD sg13g2_lv_pmos ad=0.1563p pd=1.22u as=0.147p ps=1.54u w=0.42u l=0.13u
N30 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N31 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N32 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N33 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N34 a_16048_13942# sg13g2_inv_1_0.Y a_16108_14037# VDD sg13g2_lv_pmos ad=79.8f pd=0.8u as=0.204p ps=1.835u w=0.42u l=0.13u
N35 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N36 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N37 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N38 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N39 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N40 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N41 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N42 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N43 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N44 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N45 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N46 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N47 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N48 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N49 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N50 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N51 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N52 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N53 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N54 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N55 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N56 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N57 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N58 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N59 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N60 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N61 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N62 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N63 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N64 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N65 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N66 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N67 a_13297_14486# a_12837_14495# a_12939_14495# VDD sg13g2_lv_pmos ad=0.41165p pd=2.12u as=0.3864p ps=2.93u w=1.12u l=0.13u
N68 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N69 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N70 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N71 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N72 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N73 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N74 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N75 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N76 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N77 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N78 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N79 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N80 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N81 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N82 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N83 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N84 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N85 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N86 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N87 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N88 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N89 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N90 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N91 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N92 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N93 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N94 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N95 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N96 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N97 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N98 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N99 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N100 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N101 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N102 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N103 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N104 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N105 sg13g2_inv_2_1.A a_17800_15272# VDD VDD sg13g2_lv_pmos ad=0.42p pd=2.99u as=0.2114p ps=1.54u w=1.12u l=0.13u
N106 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N107 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N108 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N109 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N110 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N111 a_14340_13722# sg13g2_and2_1_0.X a_14246_13722# VSS sg13g2_lv_nmos ad=60.89999f pd=0.71u as=0.1428p ps=1.52u w=0.42u l=0.13u
N112 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N113 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N114 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N115 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N116 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N117 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N118 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N119 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N120 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N121 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N122 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N123 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N124 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N125 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N126 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N127 a_15217_16349# a_14757_16007# a_14859_16007# VSS sg13g2_lv_nmos ad=0.31732p pd=1.805u as=0.2516p ps=2.16u w=0.74u l=0.13u
N128 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N129 VSS adc_done a_17800_15272# VSS sg13g2_lv_nmos ad=0.14875p pd=1.16u as=0.187p ps=1.78u w=0.55u l=0.13u
N130 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N131 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N132 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N133 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N134 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N135 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N136 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N137 a_12708_14909# a_12420_14488# a_12646_14909# VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=37.8f ps=0.6u w=0.42u l=0.13u
N138 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N139 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N140 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N141 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N142 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N143 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N144 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N145 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N146 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N147 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N148 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N149 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N150 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N151 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N152 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N153 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N154 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N155 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N156 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N157 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N158 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N159 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N160 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N161 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N162 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N163 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N164 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N165 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N166 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N167 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N168 a_14340_16000# a_14314_15964# VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0.36237p ps=2.605u w=1u l=0.13u
N169 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N170 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N171 sg13g2_buf_1_5.X a_14152_10736# VSS VSS sg13g2_lv_nmos ad=0.2886p pd=2.26u as=0.14875p ps=1.16u w=0.74u l=0.13u
N172 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N173 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N174 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N175 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N176 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N177 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N178 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N179 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N180 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N181 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N182 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N183 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N184 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N185 sg13g2_a21oi_1_0.A1 a_14538_17044# VSS VSS sg13g2_lv_nmos ad=0.2516p pd=2.16u as=0.1406p ps=1.12u w=0.74u l=0.13u
N186 sg13g2_inv_1_1.A sg13g2_a22oi_1_0.B2 a_16735_16388# VSS sg13g2_lv_nmos ad=0.2664p pd=1.46u as=0.13875p ps=1.115u w=0.74u l=0.13u
N187 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N188 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N189 sg13g2_dfrbpq_1_0.CLK a_7816_15996# VDD VDD sg13g2_lv_pmos ad=0.42p pd=2.99u as=0.2114p ps=1.54u w=1.12u l=0.13u
N190 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N191 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N192 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N193 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N194 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N195 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N196 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N197 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N198 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N199 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N200 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N201 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N202 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N203 a_13936_14726# sg13g2_inv_1_0.Y a_13996_14607# VDD sg13g2_lv_pmos ad=79.8f pd=0.8u as=0.204p ps=1.835u w=0.42u l=0.13u
N204 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N205 a_14314_15964# a_14757_16007# a_14054_16434# VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0.1296p ps=1.52u w=0.42u l=0.13u
N206 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N207 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N208 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N209 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N210 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N211 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N212 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N213 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N214 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N215 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N216 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N217 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N218 sg13g2_dfrbpq_1_5.Q a_16266_15996# VDD VDD sg13g2_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
N219 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N220 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N221 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N222 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N223 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N224 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N225 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N226 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N227 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N228 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N229 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N230 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N231 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N232 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N233 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N234 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N235 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N236 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N237 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N238 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N239 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N240 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N241 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N242 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N243 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N244 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N245 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N246 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N247 a_13456_13942# sg13g2_inv_1_0.Y a_13516_14037# VDD sg13g2_lv_pmos ad=79.8f pd=0.8u as=0.204p ps=1.835u w=0.42u l=0.13u
N248 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N249 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N250 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N251 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N252 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N253 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N254 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N255 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N256 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N257 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N258 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N259 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N260 VSS sg13g2_nor2_1_0.B sg13g2_nor2_1_0.Y VSS sg13g2_lv_nmos ad=0.2516p pd=2.16u as=0.1406p ps=1.12u w=0.74u l=0.13u
N261 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N262 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N263 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N264 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N265 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N266 a_13936_14726# a_13679_14845# a_14098_14922# VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=37.8f ps=0.6u w=0.42u l=0.13u
N267 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N268 a_14188_17061# a_14128_16966# a_14073_17061# VDD sg13g2_lv_pmos ad=0.204p pd=1.835u as=93.45f ps=0.865u w=0.42u l=0.13u
N269 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N270 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N271 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N272 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N273 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N274 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N275 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N276 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N277 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N278 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N279 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N280 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N281 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N282 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N283 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N284 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N285 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N286 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N287 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N288 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N289 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N290 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N291 a_14628_16421# a_14340_16000# a_14566_16421# VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=37.8f ps=0.6u w=0.42u l=0.13u
N292 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N293 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N294 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N295 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N296 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N297 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N298 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N299 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N300 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N301 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N302 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N303 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N304 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N305 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N306 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N307 adc_start a_17128_13760# VDD VDD sg13g2_lv_pmos ad=0.42p pd=2.99u as=0.2114p ps=1.54u w=1.12u l=0.13u
N308 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N309 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N310 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N311 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N312 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N313 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N314 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N315 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N316 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N317 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N318 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N319 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N320 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N321 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N322 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N323 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N324 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N325 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N326 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N327 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N328 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N329 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N330 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N331 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N332 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N333 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N334 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N335 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N336 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N337 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N338 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N339 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N340 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N341 a_11748_13722# sg13g2_a21o_1_0.X a_11654_13722# VSS sg13g2_lv_nmos ad=60.89999f pd=0.71u as=0.1428p ps=1.52u w=0.42u l=0.13u
N342 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N343 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N344 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N345 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N346 a_12612_17064# a_12586_16969# VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0.36237p ps=2.605u w=1u l=0.13u
N347 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N348 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N349 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N350 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N351 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N352 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N353 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N354 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N355 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N356 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N357 a_12646_14909# sg13g2_inv_1_0.Y VSS VSS sg13g2_lv_nmos ad=37.8f pd=0.6u as=0.1701p ps=1.65u w=0.42u l=0.13u
N358 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N359 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N360 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N361 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N362 a_12297_14113# a_11940_14040# VDD VDD sg13g2_lv_pmos ad=63f pd=0.72u as=0.1563p ps=1.22u w=0.42u l=0.13u
N363 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N364 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N365 a_13702_12532# sg13g2_buf_1_0.A a_13459_12404# VDD sg13g2_lv_pmos ad=0.2125p pd=1.425u as=0.35p ps=2.7u w=1u l=0.13u
N366 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N367 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N368 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N369 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N370 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N371 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N372 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N373 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N374 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N375 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N376 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N377 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N378 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N379 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N380 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N381 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N382 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N383 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N384 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N385 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N386 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N387 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N388 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N389 a_15409_14018# a_14949_13701# a_15051_13844# VDD sg13g2_lv_pmos ad=0.41165p pd=2.12u as=0.3864p ps=2.93u w=1.12u l=0.13u
N390 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N391 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N392 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N393 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N394 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N395 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N396 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N397 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N398 adc_en a_13576_4688# VSS VSS sg13g2_lv_nmos ad=0.2886p pd=2.26u as=0.14875p ps=1.16u w=0.74u l=0.13u
N399 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N400 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N401 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N402 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N403 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N404 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N405 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N406 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N407 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N408 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N409 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N410 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N411 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N412 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N413 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N414 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N415 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N416 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N417 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N418 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N419 VDD reset a_8968_13760# VDD sg13g2_lv_pmos ad=0.2114p pd=1.54u as=0.2856p ps=2.36u w=0.84u l=0.13u
N420 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N421 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N422 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N423 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N424 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N425 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N426 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N427 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N428 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N429 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N430 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N431 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N432 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N433 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N434 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N435 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N436 VDD a_15791_15311# a_16048_15454# VDD sg13g2_lv_pmos ad=0.4659p pd=3.65u as=79.8f ps=0.8u w=0.42u l=0.13u
N437 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N438 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N439 VSS a_15599_16357# a_16266_15996# VSS sg13g2_lv_nmos ad=0.1406p pd=1.12u as=0.2516p ps=2.16u w=0.74u l=0.13u
N440 sg13g2_inv_1_0.Y sg13g2_buf_1_6.X VSS VSS sg13g2_lv_nmos ad=0.2516p pd=2.16u as=0.2516p ps=2.16u w=0.74u l=0.13u
N441 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N442 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N443 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N444 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N445 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N446 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N447 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N448 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N449 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N450 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N451 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N452 clk_gating_en a_14632_4688# VDD VDD sg13g2_lv_pmos ad=0.42p pd=2.99u as=0.2114p ps=1.54u w=1.12u l=0.13u
N453 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N454 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N455 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N456 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N457 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N458 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N459 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N460 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N461 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N462 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N463 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N464 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N465 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N466 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N467 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N468 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N469 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N470 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N471 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N472 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N473 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N474 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N475 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N476 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N477 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N478 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N479 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N480 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N481 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N482 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N483 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N484 a_11493_16007# sg13g2_dfrbpq_1_0.CLK a_11953_16349# VSS sg13g2_lv_nmos ad=0.2516p pd=2.16u as=0.31732p ps=1.805u w=0.74u l=0.13u
N485 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N486 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N487 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N488 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N489 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N490 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N491 a_12420_14488# a_12394_14452# VSS VSS sg13g2_lv_nmos ad=0.2516p pd=2.16u as=0.1626p ps=1.415u w=0.74u l=0.13u
N492 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N493 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N494 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N495 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N496 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N497 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N498 uart_en a_14248_4688# VSS VSS sg13g2_lv_nmos ad=0.2886p pd=2.26u as=0.14875p ps=1.16u w=0.74u l=0.13u
N499 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N500 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N501 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N502 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N503 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N504 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N505 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N506 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N507 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N508 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N509 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N510 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N511 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N512 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N513 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N514 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N515 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N516 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N517 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N518 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N519 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N520 a_14340_16000# a_14859_16007# a_15599_16357# VSS sg13g2_lv_nmos ad=0.3473p pd=2.71u as=0.12665p ps=1.145u w=0.74u l=0.13u
N521 VDD a_15791_13799# a_16458_14020# VDD sg13g2_lv_pmos ad=0.2128p pd=1.5u as=0.3864p ps=2.93u w=1.12u l=0.13u
N522 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N523 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N524 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N525 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N526 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N527 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N528 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N529 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N530 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N531 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N532 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N533 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N534 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N535 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N536 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N537 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N538 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N539 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N540 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N541 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N542 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N543 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N544 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N545 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N546 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N547 a_14532_15552# a_14506_15457# VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0.36237p ps=2.605u w=1u l=0.13u
N548 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N549 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N550 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N551 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N552 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N553 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N554 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N555 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N556 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N557 a_14889_14113# a_14532_14040# VDD VDD sg13g2_lv_pmos ad=63f pd=0.72u as=0.1563p ps=1.22u w=0.42u l=0.13u
N558 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N559 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N560 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N561 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N562 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N563 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N564 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N565 VSS a_12592_16238# a_12241_16357# VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
N566 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N567 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N568 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N569 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N570 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N571 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N572 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N573 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N574 a_14073_17061# a_13131_16868# a_13871_16823# VDD sg13g2_lv_pmos ad=93.45f pd=0.865u as=0.2048p ps=1.63u w=0.42u l=0.13u
N575 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N576 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N577 a_12586_16969# a_13029_16725# a_12326_16746# VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0.1296p ps=1.52u w=0.42u l=0.13u
N578 a_12592_16238# a_12335_16357# a_12754_16434# VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=37.8f ps=0.6u w=0.42u l=0.13u
N579 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N580 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N581 VSS a_16048_13942# a_15697_13799# VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
N582 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N583 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N584 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N585 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N586 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N587 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N588 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N589 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N590 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N591 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N592 a_11433_16043# a_11076_16000# VDD VDD sg13g2_lv_pmos ad=63f pd=0.72u as=0.1563p ps=1.22u w=0.42u l=0.13u
N593 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N594 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N595 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N596 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N597 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N598 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N599 a_12817_14018# a_12357_13701# a_12459_13844# VDD sg13g2_lv_pmos ad=0.41165p pd=2.12u as=0.3864p ps=2.93u w=1.12u l=0.13u
N600 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N601 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N602 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N603 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N604 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N605 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N606 a_14532_15552# a_14506_15457# VSS VSS sg13g2_lv_nmos ad=0.2516p pd=2.16u as=0.1626p ps=1.415u w=0.74u l=0.13u
N607 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N608 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N609 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N610 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N611 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N612 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N613 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N614 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N615 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N616 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N617 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N618 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N619 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N620 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N621 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N622 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N623 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N624 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N625 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N626 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N627 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N628 a_13679_14845# a_12837_14495# a_13585_14845# VSS sg13g2_lv_nmos ad=0.12665p pd=1.145u as=0.1428p ps=1.52u w=0.42u l=0.13u
N629 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N630 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N631 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N632 a_11050_15964# a_11493_16007# a_11433_16043# VDD sg13g2_lv_pmos ad=79.8f pd=0.8u as=63f ps=0.72u w=0.42u l=0.13u
N633 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N634 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N635 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N636 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N637 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N638 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N639 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N640 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N641 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N642 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N643 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N644 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N645 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N646 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N647 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N648 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N649 a_16735_15972# sg13g2_dfrbpq_1_3.Q VDD VDD sg13g2_lv_pmos ad=0.2716p pd=1.605u as=0.3808p ps=2.92u w=1.12u l=0.13u
N650 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N651 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N652 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N653 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N654 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N655 sg13g2_and2_1_0.X a_14061_12256# VDD VDD sg13g2_lv_pmos ad=0.3808p pd=2.92u as=0.1918p ps=1.5u w=1.12u l=0.13u
N656 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N657 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N658 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N659 a_15409_15255# a_14949_15213# a_15051_15356# VSS sg13g2_lv_nmos ad=0.31732p pd=1.805u as=0.2516p ps=2.16u w=0.74u l=0.13u
N660 a_16051_14746# sg13g2_dfrbpq_1_1.Q VSS VSS sg13g2_lv_nmos ad=0.1216p pd=1.02u as=0.15745p ps=1.175u w=0.64u l=0.13u
N661 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N662 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N663 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N664 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N665 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N666 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N667 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N668 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N669 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N670 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N671 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N672 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N673 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N674 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N675 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N676 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N677 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N678 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N679 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N680 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N681 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N682 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N683 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N684 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N685 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N686 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N687 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N688 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N689 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N690 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N691 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N692 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N693 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N694 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N695 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N696 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N697 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N698 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N699 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N700 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N701 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N702 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N703 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N704 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N705 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N706 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N707 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N708 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N709 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N710 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N711 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N712 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N713 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N714 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N715 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N716 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N717 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N718 a_15409_15530# a_14949_15213# a_15051_15356# VDD sg13g2_lv_pmos ad=0.41165p pd=2.12u as=0.3864p ps=2.93u w=1.12u l=0.13u
N719 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N720 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N721 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N722 VDD a_13199_13799# a_13866_14020# VDD sg13g2_lv_pmos ad=0.2128p pd=1.5u as=0.3864p ps=2.93u w=1.12u l=0.13u
N723 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N724 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N725 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N726 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N727 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N728 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N729 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N730 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N731 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N732 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N733 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N734 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N735 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N736 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N737 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N738 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N739 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N740 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N741 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N742 sg13g2_o21ai_1_0.B1 a_14235_17564# a_14437_17878# VSS sg13g2_lv_nmos ad=0.333p pd=2.38u as=0.1406p ps=1.12u w=0.74u l=0.13u
N743 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N744 a_12394_14452# a_12837_14495# a_12777_14531# VDD sg13g2_lv_pmos ad=79.8f pd=0.8u as=63f ps=0.72u w=0.42u l=0.13u
N745 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N746 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N747 VDD sg13g2_inv_1_0.Y a_14246_13722# VDD sg13g2_lv_pmos ad=0.36237p pd=2.605u as=79.8f ps=0.8u w=0.42u l=0.13u
N748 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N749 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N750 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N751 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N752 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N753 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N754 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N755 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N756 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N757 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N758 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N759 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N760 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N761 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N762 sc_en a_14440_5412# VSS VSS sg13g2_lv_nmos ad=0.2886p pd=2.26u as=0.14875p ps=1.16u w=0.74u l=0.13u
N763 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N764 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N765 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N766 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N767 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N768 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N769 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N770 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N771 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N772 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N773 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N774 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N775 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N776 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N777 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N778 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N779 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N780 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N781 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N782 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N783 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N784 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N785 a_13838_12256# sg13g2_buf_1_4.A a_13459_12404# VSS sg13g2_lv_nmos ad=81.6f pd=0.895u as=0.1216p ps=1.02u w=0.64u l=0.13u
N786 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N787 VDD a_13871_16823# a_14538_17044# VDD sg13g2_lv_pmos ad=0.2128p pd=1.5u as=0.3864p ps=2.93u w=1.12u l=0.13u
N788 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N789 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N790 VSS sg13g2_inv_1_0.Y a_12228_14922# VSS sg13g2_lv_nmos ad=0.1626p pd=1.415u as=60.89999f ps=0.71u w=0.42u l=0.13u
N791 VSS a_13456_13942# a_13105_13799# VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
N792 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N793 a_12900_16759# a_13131_16868# a_12586_16969# VSS sg13g2_lv_nmos ad=0.2373p pd=1.97u as=79.8f ps=0.8u w=0.42u l=0.13u
N794 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N795 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N796 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N797 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N798 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N799 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N800 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N801 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N802 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N803 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N804 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N805 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N806 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N807 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N808 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N809 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N810 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N811 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N812 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N813 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N814 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N815 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N816 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N817 a_14820_15247# a_15051_15356# a_14506_15457# VSS sg13g2_lv_nmos ad=0.2373p pd=1.97u as=79.8f ps=0.8u w=0.42u l=0.13u
N818 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N819 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N820 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N821 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N822 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N823 sg13g2_o21ai_1_0.A1 sg13g2_dfrbpq_1_5.Q VDD VDD sg13g2_lv_pmos ad=0.3808p pd=2.92u as=0.3808p ps=2.92u w=1.12u l=0.13u
N824 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N825 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N826 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N827 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N828 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N829 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N830 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N831 a_12969_17137# a_12612_17064# VDD VDD sg13g2_lv_pmos ad=63f pd=0.72u as=0.1563p ps=1.22u w=0.42u l=0.13u
N832 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N833 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N834 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N835 VSS reset a_8968_13760# VSS sg13g2_lv_nmos ad=0.14875p pd=1.16u as=0.187p ps=1.78u w=0.55u l=0.13u
N836 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N837 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N838 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N839 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N840 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N841 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N842 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N843 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N844 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N845 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N846 adc_en a_13576_4688# VDD VDD sg13g2_lv_pmos ad=0.42p pd=2.99u as=0.2114p ps=1.54u w=1.12u l=0.13u
N847 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N848 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N849 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N850 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N851 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N852 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N853 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N854 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N855 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N856 VSS timer_done a_14152_10736# VSS sg13g2_lv_nmos ad=0.14875p pd=1.16u as=0.187p ps=1.78u w=0.55u l=0.13u
N857 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N858 VSS a_14128_16966# a_13777_16823# VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
N859 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N860 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N861 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N862 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N863 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N864 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N865 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N866 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N867 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N868 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N869 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N870 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N871 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N872 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N873 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N874 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N875 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N876 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N877 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N878 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N879 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N880 sg13g2_nor2b_1_0.Y a_12046_15276# VSS VSS sg13g2_lv_nmos ad=0.1406p pd=1.12u as=0.17255p ps=1.25u w=0.74u l=0.13u
N881 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N882 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N883 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N884 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N885 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N886 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N887 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N888 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N889 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N890 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N891 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N892 sg13g2_dfrbpq_1_3.Q a_16458_15532# VDD VDD sg13g2_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
N893 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N894 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N895 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N896 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N897 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N898 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N899 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N900 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N901 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N902 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N903 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N904 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N905 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N906 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N907 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N908 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N909 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N910 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N911 a_12420_14488# a_12394_14452# VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0.36237p ps=2.605u w=1u l=0.13u
N912 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N913 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N914 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N915 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N916 a_12537_16119# a_11595_16007# a_12335_16357# VDD sg13g2_lv_pmos ad=93.45f pd=0.865u as=0.2048p ps=1.63u w=0.42u l=0.13u
N917 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N918 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N919 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N920 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N921 sg13g2_inv_1_0.Y sg13g2_buf_1_6.X VDD VDD sg13g2_lv_pmos ad=0.3808p pd=2.92u as=0.3808p ps=2.92u w=1.12u l=0.13u
N922 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N923 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N924 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N925 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N926 a_14532_15552# a_15051_15356# a_15791_15311# VSS sg13g2_lv_nmos ad=0.3473p pd=2.71u as=0.12665p ps=1.145u w=0.74u l=0.13u
N927 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N928 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N929 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N930 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N931 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N932 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N933 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N934 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N935 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N936 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N937 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N938 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N939 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N940 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N941 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N942 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N943 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N944 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N945 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N946 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N947 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N948 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N949 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N950 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N951 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N952 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N953 uart_en a_14248_4688# VDD VDD sg13g2_lv_pmos ad=0.42p pd=2.99u as=0.2114p ps=1.54u w=1.12u l=0.13u
N954 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N955 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N956 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N957 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N958 sg13g2_a21o_1_0.A2 sg13g2_buf_1_5.X VSS VSS sg13g2_lv_nmos ad=0.1406p pd=1.12u as=0.2516p ps=2.16u w=0.74u l=0.13u
N959 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N960 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N961 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N962 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N963 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N964 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N965 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N966 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N967 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N968 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N969 VDD sg13g2_inv_1_0.Y a_11654_13722# VDD sg13g2_lv_pmos ad=0.36237p pd=2.605u as=79.8f ps=0.8u w=0.42u l=0.13u
N970 a_17006_16388# sg13g2_dfrbpq_1_3.Q sg13g2_inv_1_1.A VSS sg13g2_lv_nmos ad=96.2f pd=1u as=0.2664p ps=1.46u w=0.74u l=0.13u
N971 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N972 a_15791_15311# a_14949_15213# a_15697_15311# VSS sg13g2_lv_nmos ad=0.12665p pd=1.145u as=0.1428p ps=1.52u w=0.42u l=0.13u
N973 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N974 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N975 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N976 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N977 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N978 a_15916_16119# a_15856_16238# a_15801_16119# VDD sg13g2_lv_pmos ad=0.204p pd=1.835u as=93.45f ps=0.865u w=0.42u l=0.13u
N979 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N980 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N981 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N982 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N983 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N984 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N985 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N986 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N987 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N988 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N989 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N990 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N991 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N992 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N993 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N994 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N995 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N996 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N997 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N998 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N999 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1000 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1001 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1002 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1003 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1004 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1005 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1006 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1007 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1008 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1009 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1010 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1011 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1012 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1013 VDD sg13g2_buf_1_0.A a_14632_4688# VDD sg13g2_lv_pmos ad=0.2114p pd=1.54u as=0.2856p ps=2.36u w=0.84u l=0.13u
N1014 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1015 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1016 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1017 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1018 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1019 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1020 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1021 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1022 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1023 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1024 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1025 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1026 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1027 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1028 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1029 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1030 sg13g2_buf_1_6.X a_8968_13760# VDD VDD sg13g2_lv_pmos ad=0.42p pd=2.99u as=0.2114p ps=1.54u w=1.12u l=0.13u
N1031 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1032 a_14506_15457# a_14949_15213# a_14246_15234# VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0.1296p ps=1.52u w=0.42u l=0.13u
N1033 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1034 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1035 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1036 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1037 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1038 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1039 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1040 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1041 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1042 a_14820_15247# a_14532_15552# a_14758_15247# VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=37.8f ps=0.6u w=0.42u l=0.13u
N1043 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1044 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1045 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1046 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1047 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1048 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1049 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1050 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1051 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1052 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1053 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1054 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1055 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1056 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1057 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1058 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1059 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1060 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1061 VSS uart_done a_13960_25068# VSS sg13g2_lv_nmos ad=0.14875p pd=1.16u as=0.187p ps=1.78u w=0.55u l=0.13u
N1062 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1063 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1064 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1065 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1066 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1067 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1068 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1069 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1070 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1071 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1072 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1073 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1074 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1075 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1076 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1077 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1078 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1079 VSS sg13g2_inv_1_0.Y a_11748_13722# VSS sg13g2_lv_nmos ad=0.1626p pd=1.415u as=60.89999f ps=0.71u w=0.42u l=0.13u
N1080 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1081 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1082 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1083 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1084 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1085 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1086 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1087 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1088 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1089 a_11076_16000# a_11595_16007# a_12335_16357# VSS sg13g2_lv_nmos ad=0.3473p pd=2.71u as=0.12665p ps=1.145u w=0.74u l=0.13u
N1090 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1091 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1092 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1093 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1094 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1095 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1096 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1097 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1098 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1099 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1100 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1101 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1102 a_12837_14495# sg13g2_dfrbpq_1_0.CLK a_13297_14486# VDD sg13g2_lv_pmos ad=0.4088p pd=2.97u as=0.41165p ps=2.12u w=1.12u l=0.13u
N1103 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1104 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1105 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1106 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1107 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1108 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1109 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1110 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1111 VDD sg13g2_inv_1_0.Y a_12586_16969# VDD sg13g2_lv_pmos ad=0.1563p pd=1.22u as=0.147p ps=1.54u w=0.42u l=0.13u
N1112 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1113 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1114 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1115 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1116 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1117 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1118 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1119 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1120 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1121 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1122 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1123 sg13g2_a22oi_1_0.B2 a_15976_25068# VDD VDD sg13g2_lv_pmos ad=0.42p pd=2.99u as=0.2114p ps=1.54u w=1.12u l=0.13u
N1124 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1125 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1126 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1127 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1128 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1129 VDD a_14235_17564# sg13g2_o21ai_1_0.B1 VDD sg13g2_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
N1130 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1131 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1132 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1133 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1134 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1135 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1136 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1137 a_11953_16349# a_11493_16007# a_11595_16007# VSS sg13g2_lv_nmos ad=0.31732p pd=1.805u as=0.2516p ps=2.16u w=0.74u l=0.13u
N1138 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1139 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1140 a_12268_15532# a_12046_15276# VDD VDD sg13g2_lv_pmos ad=0.1176p pd=1.33u as=0.2618p ps=1.63u w=1.12u l=0.13u
N1141 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1142 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1143 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1144 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1145 a_13199_13799# a_12357_13701# a_13105_13799# VSS sg13g2_lv_nmos ad=0.12665p pd=1.145u as=0.1428p ps=1.52u w=0.42u l=0.13u
N1146 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1147 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1148 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1149 a_13601_16344# sg13g2_a21oi_1_0.A1 sg13g2_dfrbpq_1_4.D VSS sg13g2_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
N1150 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1151 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1152 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1153 a_16018_16434# sg13g2_inv_1_0.Y VSS VSS sg13g2_lv_nmos ad=37.8f pd=0.6u as=79.8f ps=0.8u w=0.42u l=0.13u
N1154 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1155 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1156 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1157 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1158 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1159 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1160 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1161 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1162 a_14757_16007# sg13g2_dfrbpq_1_0.CLK a_15217_16349# VSS sg13g2_lv_nmos ad=0.2516p pd=2.16u as=0.31732p ps=1.805u w=0.74u l=0.13u
N1163 a_16210_15234# sg13g2_inv_1_0.Y VSS VSS sg13g2_lv_nmos ad=37.8f pd=0.6u as=79.8f ps=0.8u w=0.42u l=0.13u
N1164 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1165 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1166 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1167 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1168 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1169 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1170 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1171 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1172 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1173 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1174 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1175 VDD a_12335_16357# a_13002_15996# VDD sg13g2_lv_pmos ad=0.2128p pd=1.5u as=0.3864p ps=2.93u w=1.12u l=0.13u
N1176 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1177 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1178 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1179 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1180 VDD sg13g2_inv_1_0.Y a_14054_16434# VDD sg13g2_lv_pmos ad=0.36237p pd=2.605u as=79.8f ps=0.8u w=0.42u l=0.13u
N1181 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1182 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1183 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1184 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1185 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1186 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1187 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1188 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1189 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1190 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1191 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1192 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1193 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1194 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1195 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1196 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1197 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1198 a_14532_14040# a_14506_13945# VSS VSS sg13g2_lv_nmos ad=0.2516p pd=2.16u as=0.1626p ps=1.415u w=0.74u l=0.13u
N1199 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1200 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1201 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1202 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1203 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1204 VSS a_16051_14746# sg13g2_dfrbpq_1_3.D VSS sg13g2_lv_nmos ad=0.15745p pd=1.175u as=0.2351p ps=2.16u w=0.74u l=0.13u
N1205 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1206 VDD a_15791_13799# a_16048_13942# VDD sg13g2_lv_pmos ad=0.4659p pd=3.65u as=79.8f ps=0.8u w=0.42u l=0.13u
N1207 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1208 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1209 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1210 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1211 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1212 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1213 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1214 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1215 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1216 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1217 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1218 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1219 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1220 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1221 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1222 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1223 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1224 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1225 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1226 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1227 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1228 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1229 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1230 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1231 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1232 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1233 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1234 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1235 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1236 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1237 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1238 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1239 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1240 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1241 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1242 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1243 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1244 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1245 VSS sg13g2_buf_1_0.A a_14632_4688# VSS sg13g2_lv_nmos ad=0.14875p pd=1.16u as=0.187p ps=1.78u w=0.55u l=0.13u
N1246 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1247 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1248 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1249 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1250 a_15409_13743# a_14949_13701# a_15051_13844# VSS sg13g2_lv_nmos ad=0.31732p pd=1.805u as=0.2516p ps=2.16u w=0.74u l=0.13u
N1251 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1252 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1253 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1254 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1255 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1256 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1257 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1258 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1259 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1260 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1261 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1262 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1263 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1264 a_14758_15247# sg13g2_inv_1_0.Y VSS VSS sg13g2_lv_nmos ad=37.8f pd=0.6u as=0.1701p ps=1.65u w=0.42u l=0.13u
N1265 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1266 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1267 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1268 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1269 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1270 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1271 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1272 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1273 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1274 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1275 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1276 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1277 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1278 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1279 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1280 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1281 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1282 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1283 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1284 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1285 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1286 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1287 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1288 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1289 a_15801_16119# a_14859_16007# a_15599_16357# VDD sg13g2_lv_pmos ad=93.45f pd=0.865u as=0.2048p ps=1.63u w=0.42u l=0.13u
N1290 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1291 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1292 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1293 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1294 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1295 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1296 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1297 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1298 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1299 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1300 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1301 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1302 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1303 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1304 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1305 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1306 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1307 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1308 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1309 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1310 a_11076_16000# a_11050_15964# VSS VSS sg13g2_lv_nmos ad=0.2516p pd=2.16u as=0.1626p ps=1.415u w=0.74u l=0.13u
N1311 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1312 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1313 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1314 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1315 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1316 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1317 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1318 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1319 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1320 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1321 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1322 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1323 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1324 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1325 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1326 a_11940_14040# a_12459_13844# a_13199_13799# VSS sg13g2_lv_nmos ad=0.3473p pd=2.71u as=0.12665p ps=1.145u w=0.74u l=0.13u
N1327 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1328 VDD sg13g2_inv_1_0.Y a_14506_15457# VDD sg13g2_lv_pmos ad=0.1563p pd=1.22u as=0.147p ps=1.54u w=0.42u l=0.13u
N1329 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1330 a_14532_14040# a_14506_13945# VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0.36237p ps=2.605u w=1u l=0.13u
N1331 a_13499_15996# sg13g2_nor2_1_0.Y sg13g2_dfrbpq_1_4.D VDD sg13g2_lv_pmos ad=0.2128p pd=1.5u as=0.3808p ps=2.92u w=1.12u l=0.13u
N1332 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1333 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1334 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1335 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1336 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1337 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1338 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1339 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1340 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1341 a_12228_14922# sg13g2_nor2b_1_0.Y a_12134_14922# VSS sg13g2_lv_nmos ad=60.89999f pd=0.71u as=0.1428p ps=1.52u w=0.42u l=0.13u
N1342 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1343 a_12612_17064# a_12586_16969# VSS VSS sg13g2_lv_nmos ad=0.2516p pd=2.16u as=0.1626p ps=1.415u w=0.74u l=0.13u
N1344 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1345 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1346 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1347 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1348 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1349 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1350 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1351 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1352 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1353 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1354 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1355 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1356 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1357 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1358 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1359 tx_start a_14248_23556# VDD VDD sg13g2_lv_pmos ad=0.42p pd=2.99u as=0.2114p ps=1.54u w=1.12u l=0.13u
N1360 a_15791_13799# a_14949_13701# a_15697_13799# VSS sg13g2_lv_nmos ad=0.12665p pd=1.145u as=0.1428p ps=1.52u w=0.42u l=0.13u
N1361 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1362 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1363 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1364 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1365 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1366 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1367 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1368 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1369 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1370 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1371 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1372 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1373 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1374 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1375 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1376 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1377 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1378 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1379 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1380 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1381 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1382 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1383 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1384 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1385 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1386 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1387 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1388 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1389 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1390 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1391 VDD a_13679_14845# a_13936_14726# VDD sg13g2_lv_pmos ad=0.4659p pd=3.65u as=79.8f ps=0.8u w=0.42u l=0.13u
N1392 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1393 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1394 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1395 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1396 a_14628_16421# a_14859_16007# a_14314_15964# VSS sg13g2_lv_nmos ad=0.2373p pd=1.97u as=79.8f ps=0.8u w=0.42u l=0.13u
N1397 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1398 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1399 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1400 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1401 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1402 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1403 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1404 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1405 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1406 a_15217_15998# a_14757_16007# a_14859_16007# VDD sg13g2_lv_pmos ad=0.41165p pd=2.12u as=0.3864p ps=2.93u w=1.12u l=0.13u
N1407 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1408 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1409 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1410 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1411 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1412 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1413 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1414 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1415 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1416 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1417 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1418 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1419 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1420 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1421 a_11914_13945# a_12357_13701# a_11654_13722# VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0.1296p ps=1.52u w=0.42u l=0.13u
N1422 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1423 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1424 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1425 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1426 a_11940_14040# a_11914_13945# VSS VSS sg13g2_lv_nmos ad=0.2516p pd=2.16u as=0.1626p ps=1.415u w=0.74u l=0.13u
N1427 a_14820_13735# a_15051_13844# a_14506_13945# VSS sg13g2_lv_nmos ad=0.2373p pd=1.97u as=79.8f ps=0.8u w=0.42u l=0.13u
N1428 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1429 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1430 a_14949_13701# sg13g2_dfrbpq_1_0.CLK a_15409_14018# VDD sg13g2_lv_pmos ad=0.4088p pd=2.97u as=0.41165p ps=2.12u w=1.12u l=0.13u
N1431 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1432 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1433 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1434 VDD a_13199_13799# a_13456_13942# VDD sg13g2_lv_pmos ad=0.4659p pd=3.65u as=79.8f ps=0.8u w=0.42u l=0.13u
N1435 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1436 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1437 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1438 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1439 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1440 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1441 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1442 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1443 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1444 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1445 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1446 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1447 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1448 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1449 VDD sg13g2_buf_1_0.A a_13576_4688# VDD sg13g2_lv_pmos ad=0.2114p pd=1.54u as=0.2856p ps=2.36u w=0.84u l=0.13u
N1450 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1451 a_14128_16966# sg13g2_inv_1_0.Y a_14188_17061# VDD sg13g2_lv_pmos ad=79.8f pd=0.8u as=0.204p ps=1.835u w=0.42u l=0.13u
N1452 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1453 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1454 VDD clk a_7816_15996# VDD sg13g2_lv_pmos ad=0.2114p pd=1.54u as=0.2856p ps=2.36u w=0.84u l=0.13u
N1455 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1456 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1457 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1458 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1459 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1460 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1461 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1462 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1463 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1464 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1465 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1466 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1467 sg13g2_o21ai_1_0.A1 sg13g2_dfrbpq_1_5.Q VSS VSS sg13g2_lv_nmos ad=0.2516p pd=2.16u as=0.2516p ps=2.16u w=0.74u l=0.13u
N1468 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1469 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1470 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1471 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1472 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1473 VSS sg13g2_inv_2_1.A a_17006_16388# VSS sg13g2_lv_nmos ad=0.2516p pd=2.16u as=96.2f ps=1u w=0.74u l=0.13u
N1474 a_12817_13743# a_12357_13701# a_12459_13844# VSS sg13g2_lv_nmos ad=0.31732p pd=1.805u as=0.2516p ps=2.16u w=0.74u l=0.13u
N1475 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1476 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1477 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1478 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1479 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1480 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1481 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1482 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1483 sg13g2_buf_1_4.A a_13866_14020# VDD VDD sg13g2_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
N1484 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1485 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1486 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1487 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1488 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1489 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1490 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1491 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1492 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1493 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1494 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1495 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1496 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1497 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1498 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1499 VDD a_13679_14845# a_14346_14484# VDD sg13g2_lv_pmos ad=0.2128p pd=1.5u as=0.3864p ps=2.93u w=1.12u l=0.13u
N1500 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1501 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1502 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1503 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1504 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1505 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1506 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1507 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1508 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1509 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1510 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1511 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1512 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1513 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1514 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1515 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1516 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1517 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1518 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1519 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1520 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1521 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1522 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1523 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1524 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1525 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1526 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1527 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1528 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1529 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1530 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1531 a_14532_14040# a_15051_13844# a_15791_13799# VSS sg13g2_lv_nmos ad=0.3473p pd=2.71u as=0.12665p ps=1.145u w=0.74u l=0.13u
N1532 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1533 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1534 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1535 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1536 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1537 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1538 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1539 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1540 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1541 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1542 VDD sg13g2_buf_1_0.A a_14248_4688# VDD sg13g2_lv_pmos ad=0.2114p pd=1.54u as=0.2856p ps=2.36u w=0.84u l=0.13u
N1543 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1544 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1545 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1546 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1547 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1548 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1549 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1550 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1551 a_13489_16767# a_13029_16725# a_13131_16868# VSS sg13g2_lv_nmos ad=0.31732p pd=1.805u as=0.2516p ps=2.16u w=0.74u l=0.13u
N1552 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1553 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1554 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1555 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1556 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1557 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1558 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1559 a_11940_14040# a_11914_13945# VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0.36237p ps=2.605u w=1u l=0.13u
N1560 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1561 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1562 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1563 VDD sg13g2_inv_1_0.Y a_14314_15964# VDD sg13g2_lv_pmos ad=0.1563p pd=1.22u as=0.147p ps=1.54u w=0.42u l=0.13u
N1564 VSS a_13679_14845# a_14346_14484# VSS sg13g2_lv_nmos ad=0.1406p pd=1.12u as=0.2516p ps=2.16u w=0.74u l=0.13u
N1565 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1566 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1567 VDD timer_done a_14152_10736# VDD sg13g2_lv_pmos ad=0.2114p pd=1.54u as=0.2856p ps=2.36u w=0.84u l=0.13u
N1568 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1569 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1570 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1571 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1572 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1573 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1574 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1575 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1576 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1577 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1578 sg13g2_dfrbpq_1_0.CLK a_7816_15996# VSS VSS sg13g2_lv_nmos ad=0.2886p pd=2.26u as=0.14875p ps=1.16u w=0.74u l=0.13u
N1579 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1580 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1581 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1582 a_12652_16119# a_12592_16238# a_12537_16119# VDD sg13g2_lv_pmos ad=0.204p pd=1.835u as=93.45f ps=0.865u w=0.42u l=0.13u
N1583 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1584 VSS sg13g2_a21o_1_0.A2 a_13838_12256# VSS sg13g2_lv_nmos ad=0.2176p pd=1.96u as=81.6f ps=0.895u w=0.64u l=0.13u
N1585 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1586 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1587 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1588 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1589 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1590 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1591 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1592 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1593 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1594 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1595 a_16294_14484# sg13g2_dfrbpq_1_1.Q a_16051_14746# VDD sg13g2_lv_pmos ad=0.2125p pd=1.425u as=0.35p ps=2.7u w=1u l=0.13u
N1596 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1597 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1598 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1599 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1600 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1601 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1602 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1603 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1604 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1605 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1606 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1607 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1608 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1609 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1610 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1611 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1612 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1613 sg13g2_dfrbpq_1_5.Q a_16266_15996# VSS VSS sg13g2_lv_nmos ad=0.2516p pd=2.16u as=0.1406p ps=1.12u w=0.74u l=0.13u
N1614 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1615 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1616 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1617 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1618 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1619 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1620 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1621 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1622 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1623 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1624 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1625 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1626 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1627 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1628 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1629 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1630 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1631 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1632 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1633 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1634 a_14506_13945# a_14949_13701# a_14246_13722# VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0.1296p ps=1.52u w=0.42u l=0.13u
N1635 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1636 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1637 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1638 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1639 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1640 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1641 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1642 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1643 a_14820_13735# a_14532_14040# a_14758_13735# VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=37.8f ps=0.6u w=0.42u l=0.13u
N1644 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1645 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1646 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1647 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1648 a_12166_13735# sg13g2_inv_1_0.Y VSS VSS sg13g2_lv_nmos ad=37.8f pd=0.6u as=0.1701p ps=1.65u w=0.42u l=0.13u
N1649 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1650 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1651 a_12357_13701# sg13g2_dfrbpq_1_0.CLK a_12817_14018# VDD sg13g2_lv_pmos ad=0.4088p pd=2.97u as=0.41165p ps=2.12u w=1.12u l=0.13u
N1652 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1653 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1654 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1655 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1656 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1657 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1658 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1659 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1660 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1661 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1662 VSS sg13g2_a21o_1_1.A2 a_16430_14832# VSS sg13g2_lv_nmos ad=0.2176p pd=1.96u as=81.6f ps=0.895u w=0.64u l=0.13u
N1663 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1664 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1665 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1666 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1667 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1668 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1669 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1670 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1671 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1672 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1673 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1674 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1675 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1676 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1677 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1678 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1679 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1680 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1681 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1682 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1683 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1684 VSS sg13g2_buf_1_0.A a_13576_4688# VSS sg13g2_lv_nmos ad=0.14875p pd=1.16u as=0.187p ps=1.78u w=0.55u l=0.13u
N1685 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1686 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1687 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1688 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1689 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1690 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1691 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1692 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1693 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1694 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1695 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1696 sg13g2_dfrbpq_1_1.Q a_16458_14020# VDD VDD sg13g2_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
N1697 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1698 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1699 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1700 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1701 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1702 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1703 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1704 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1705 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1706 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1707 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1708 sg13g2_inv_1_1.A sg13g2_dfrbpq_1_5.Q a_16735_15972# VDD sg13g2_lv_pmos ad=0.2128p pd=1.5u as=0.2716p ps=1.605u w=1.12u l=0.13u
N1709 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1710 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1711 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1712 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1713 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1714 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1715 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1716 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1717 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1718 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1719 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1720 a_14949_15213# sg13g2_dfrbpq_1_0.CLK a_15409_15255# VSS sg13g2_lv_nmos ad=0.2516p pd=2.16u as=0.31732p ps=1.805u w=0.74u l=0.13u
N1721 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1722 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1723 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1724 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1725 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1726 VSS sg13g2_buf_1_5.X sg13g2_a21o_1_0.A2 VSS sg13g2_lv_nmos ad=0.2516p pd=2.16u as=0.1406p ps=1.12u w=0.74u l=0.13u
N1727 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1728 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1729 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1730 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1731 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1732 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1733 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1734 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1735 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1736 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1737 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1738 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1739 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1740 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1741 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1742 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1743 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1744 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1745 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1746 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1747 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1748 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1749 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1750 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1751 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1752 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1753 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1754 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1755 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1756 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1757 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1758 a_12754_16434# sg13g2_inv_1_0.Y VSS VSS sg13g2_lv_nmos ad=37.8f pd=0.6u as=79.8f ps=0.8u w=0.42u l=0.13u
N1759 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1760 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1761 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1762 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1763 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1764 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1765 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1766 VDD sg13g2_buf_1_4.A a_13702_12532# VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0.2125p ps=1.425u w=1u l=0.13u
N1767 a_11493_16007# sg13g2_dfrbpq_1_0.CLK a_11953_15998# VDD sg13g2_lv_pmos ad=0.4088p pd=2.97u as=0.41165p ps=2.12u w=1.12u l=0.13u
N1768 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1769 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1770 a_16210_13722# sg13g2_inv_1_0.Y VSS VSS sg13g2_lv_nmos ad=37.8f pd=0.6u as=79.8f ps=0.8u w=0.42u l=0.13u
N1771 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1772 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1773 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1774 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1775 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1776 VSS sg13g2_buf_1_0.A a_14248_4688# VSS sg13g2_lv_nmos ad=0.14875p pd=1.16u as=0.187p ps=1.78u w=0.55u l=0.13u
N1777 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1778 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1779 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1780 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1781 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1782 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1783 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1784 sg13g2_buf_1_5.X a_14152_10736# VDD VDD sg13g2_lv_pmos ad=0.42p pd=2.99u as=0.2114p ps=1.54u w=1.12u l=0.13u
N1785 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1786 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1787 a_14949_15213# sg13g2_dfrbpq_1_0.CLK a_15409_15530# VDD sg13g2_lv_pmos ad=0.4088p pd=2.97u as=0.41165p ps=2.12u w=1.12u l=0.13u
N1788 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1789 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1790 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1791 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1792 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1793 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1794 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1795 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1796 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1797 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1798 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1799 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1800 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1801 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1802 sg13g2_and2_1_0.X a_14061_12256# VSS VSS sg13g2_lv_nmos ad=0.2516p pd=2.16u as=0.1331p ps=1.12u w=0.74u l=0.13u
N1803 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1804 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1805 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1806 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1807 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1808 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1809 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1810 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1811 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1812 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1813 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1814 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1815 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1816 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1817 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1818 a_13489_17042# a_13029_16725# a_13131_16868# VDD sg13g2_lv_pmos ad=0.41165p pd=2.12u as=0.3864p ps=2.93u w=1.12u l=0.13u
N1819 a_15856_16238# a_15599_16357# a_16018_16434# VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=37.8f ps=0.6u w=0.42u l=0.13u
N1820 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1821 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1822 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1823 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1824 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1825 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1826 a_10790_16434# a_11595_16007# a_11050_15964# VDD sg13g2_lv_pmos ad=0.1428p pd=1.52u as=79.8f ps=0.8u w=0.42u l=0.13u
N1827 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1828 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1829 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1830 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1831 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1832 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1833 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1834 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1835 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1836 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1837 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1838 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1839 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1840 a_12612_17064# a_13131_16868# a_13871_16823# VSS sg13g2_lv_nmos ad=0.3473p pd=2.71u as=0.12665p ps=1.145u w=0.74u l=0.13u
N1841 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1842 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1843 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1844 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1845 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1846 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1847 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1848 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1849 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1850 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1851 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1852 Timer_en a_13768_10736# VSS VSS sg13g2_lv_nmos ad=0.2886p pd=2.26u as=0.14875p ps=1.16u w=0.74u l=0.13u
N1853 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1854 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1855 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1856 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1857 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1858 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1859 a_16430_14832# sg13g2_dfrbpq_1_3.Q a_16051_14746# VSS sg13g2_lv_nmos ad=81.6f pd=0.895u as=0.1216p ps=1.02u w=0.64u l=0.13u
N1860 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1861 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1862 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1863 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1864 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1865 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1866 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1867 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1868 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1869 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1870 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1871 VDD sg13g2_buf_1_0.A a_14440_5412# VDD sg13g2_lv_pmos ad=0.2114p pd=1.54u as=0.2856p ps=2.36u w=0.84u l=0.13u
N1872 a_14155_12256# sg13g2_buf_1_4.A a_14061_12256# VSS sg13g2_lv_nmos ad=0.1216p pd=1.02u as=0.2176p ps=1.96u w=0.64u l=0.13u
N1873 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1874 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1875 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1876 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1877 a_14246_15234# a_15051_15356# a_14506_15457# VDD sg13g2_lv_pmos ad=0.1428p pd=1.52u as=79.8f ps=0.8u w=0.42u l=0.13u
N1878 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1879 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1880 a_14758_13735# sg13g2_inv_1_0.Y VSS VSS sg13g2_lv_nmos ad=37.8f pd=0.6u as=0.1701p ps=1.65u w=0.42u l=0.13u
N1881 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1882 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1883 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1884 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1885 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1886 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1887 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1888 a_16108_15549# a_16048_15454# a_15993_15549# VDD sg13g2_lv_pmos ad=0.204p pd=1.835u as=93.45f ps=0.865u w=0.42u l=0.13u
N1889 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1890 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1891 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1892 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1893 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1894 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1895 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1896 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1897 a_13871_16823# a_13029_16725# a_13777_16823# VSS sg13g2_lv_nmos ad=0.12665p pd=1.145u as=0.1428p ps=1.52u w=0.42u l=0.13u
N1898 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1899 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1900 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1901 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1902 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1903 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1904 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1905 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1906 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1907 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1908 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1909 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1910 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1911 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1912 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1913 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1914 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1915 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1916 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1917 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1918 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1919 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1920 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1921 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1922 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1923 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1924 VDD sg13g2_inv_1_0.Y a_11914_13945# VDD sg13g2_lv_pmos ad=0.1563p pd=1.22u as=0.147p ps=1.54u w=0.42u l=0.13u
N1925 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1926 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1927 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1928 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1929 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1930 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1931 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1932 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1933 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1934 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1935 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1936 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1937 VSS a_15791_15311# a_16458_15532# VSS sg13g2_lv_nmos ad=0.1406p pd=1.12u as=0.2516p ps=2.16u w=0.74u l=0.13u
N1938 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1939 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1940 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1941 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1942 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1943 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1944 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1945 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1946 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1947 a_12134_14922# a_12939_14495# a_12394_14452# VDD sg13g2_lv_pmos ad=0.1428p pd=1.52u as=79.8f ps=0.8u w=0.42u l=0.13u
N1948 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1949 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1950 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1951 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1952 a_12900_16759# a_12612_17064# a_12838_16759# VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=37.8f ps=0.6u w=0.42u l=0.13u
N1953 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1954 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1955 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1956 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1957 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1958 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1959 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1960 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1961 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1962 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1963 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1964 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1965 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1966 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1967 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1968 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1969 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1970 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1971 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1972 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1973 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1974 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1975 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1976 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1977 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1978 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1979 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1980 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1981 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1982 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1983 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1984 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1985 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1986 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1987 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1988 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1989 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1990 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1991 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N1992 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1993 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N1994 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1995 sg13g2_a21oi_1_0.A1 a_14538_17044# VDD VDD sg13g2_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
N1996 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N1997 VDD sg13g2_nor2_1_0.A a_12046_15276# VDD sg13g2_lv_pmos ad=0.2618p pd=1.63u as=0.2856p ps=2.36u w=0.84u l=0.13u
N1998 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N1999 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2000 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2001 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2002 a_13618_13722# sg13g2_inv_1_0.Y VSS VSS sg13g2_lv_nmos ad=37.8f pd=0.6u as=79.8f ps=0.8u w=0.42u l=0.13u
N2003 VDD sg13g2_a21oi_1_0.A2 a_14235_17564# VDD sg13g2_lv_pmos ad=0.2198p pd=1.53u as=0.2856p ps=2.36u w=0.84u l=0.13u
N2004 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2005 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2006 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2007 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2008 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2009 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2010 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2011 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2012 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2013 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2014 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2015 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2016 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2017 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2018 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2019 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2020 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2021 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2022 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2023 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2024 a_14340_16000# a_14314_15964# VSS VSS sg13g2_lv_nmos ad=0.2516p pd=2.16u as=0.1626p ps=1.415u w=0.74u l=0.13u
N2025 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2026 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2027 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2028 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2029 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2030 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2031 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2032 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2033 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2034 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2035 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2036 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2037 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2038 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2039 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2040 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2041 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2042 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2043 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2044 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2045 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2046 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2047 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2048 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2049 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2050 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2051 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2052 sg13g2_nor2b_1_0.Y sg13g2_nor2_1_0.B a_12268_15532# VDD sg13g2_lv_pmos ad=0.3808p pd=2.92u as=0.1176p ps=1.33u w=1.12u l=0.13u
N2053 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2054 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2055 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2056 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2057 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2058 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2059 sg13g2_a21o_1_1.A2 sg13g2_inv_2_1.A VSS VSS sg13g2_lv_nmos ad=0.1406p pd=1.12u as=0.2516p ps=2.16u w=0.74u l=0.13u
N2060 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2061 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2062 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2063 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2064 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2065 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2066 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2067 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2068 a_14506_15457# a_14949_15213# a_14889_15625# VDD sg13g2_lv_pmos ad=79.8f pd=0.8u as=63f ps=0.72u w=0.42u l=0.13u
N2069 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2070 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2071 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2072 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2073 a_14290_16746# sg13g2_inv_1_0.Y VSS VSS sg13g2_lv_nmos ad=37.8f pd=0.6u as=79.8f ps=0.8u w=0.42u l=0.13u
N2074 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2075 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2076 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2077 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2078 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2079 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2080 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2081 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2082 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2083 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2084 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2085 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2086 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2087 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2088 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2089 VSS sg13g2_nor2_1_0.B sg13g2_nor2b_1_0.Y VSS sg13g2_lv_nmos ad=0.2516p pd=2.16u as=0.1406p ps=1.12u w=0.74u l=0.13u
N2090 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2091 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2092 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2093 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2094 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2095 VSS sg13g2_buf_1_5.X a_14155_12256# VSS sg13g2_lv_nmos ad=0.1331p pd=1.12u as=0.1216p ps=1.02u w=0.64u l=0.13u
N2096 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2097 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2098 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2099 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2100 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2101 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2102 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2103 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2104 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2105 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2106 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2107 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2108 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2109 VSS sg13g2_nor2_1_0.A a_12046_15276# VSS sg13g2_lv_nmos ad=0.17255p pd=1.25u as=0.187p ps=1.78u w=0.55u l=0.13u
N2110 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2111 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2112 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2113 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2114 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2115 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2116 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2117 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2118 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2119 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2120 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2121 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2122 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2123 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2124 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2125 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2126 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2127 VDD sg13g2_inv_1_0.Y a_14506_13945# VDD sg13g2_lv_pmos ad=0.1563p pd=1.22u as=0.147p ps=1.54u w=0.42u l=0.13u
N2128 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2129 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2130 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2131 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2132 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2133 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2134 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2135 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2136 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2137 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2138 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2139 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2140 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2141 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2142 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2143 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2144 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2145 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2146 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2147 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2148 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2149 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2150 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2151 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2152 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2153 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2154 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2155 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2156 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2157 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2158 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2159 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2160 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2161 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2162 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2163 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2164 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2165 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2166 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2167 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2168 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2169 a_12838_16759# sg13g2_inv_1_0.Y VSS VSS sg13g2_lv_nmos ad=37.8f pd=0.6u as=0.1701p ps=1.65u w=0.42u l=0.13u
N2170 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2171 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2172 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2173 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2174 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2175 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2176 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2177 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2178 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2179 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2180 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2181 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2182 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2183 a_15599_16357# a_14757_16007# a_15505_16357# VSS sg13g2_lv_nmos ad=0.12665p pd=1.145u as=0.1428p ps=1.52u w=0.42u l=0.13u
N2184 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2185 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2186 a_15856_16238# sg13g2_inv_1_0.Y a_15916_16119# VDD sg13g2_lv_pmos ad=79.8f pd=0.8u as=0.204p ps=1.835u w=0.42u l=0.13u
N2187 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2188 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2189 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2190 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2191 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2192 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2193 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2194 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2195 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2196 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2197 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2198 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2199 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2200 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2201 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2202 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2203 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2204 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2205 VDD sg13g2_dfrbpq_1_1.Q a_17128_13760# VDD sg13g2_lv_pmos ad=0.2114p pd=1.54u as=0.2856p ps=2.36u w=0.84u l=0.13u
N2206 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2207 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2208 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2209 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2210 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2211 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2212 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2213 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2214 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2215 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2216 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2217 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2218 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2219 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2220 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2221 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2222 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2223 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2224 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2225 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2226 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2227 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2228 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2229 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2230 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2231 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2232 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2233 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2234 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2235 a_15791_15311# a_14949_15213# a_14532_15552# VDD sg13g2_lv_pmos ad=0.2048p pd=1.63u as=0.34p ps=2.68u w=1u l=0.13u
N2236 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2237 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2238 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2239 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2240 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2241 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2242 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2243 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2244 a_16048_15454# a_15791_15311# a_16210_15234# VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=37.8f ps=0.6u w=0.42u l=0.13u
N2245 VSS a_13936_14726# a_13585_14845# VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
N2246 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2247 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2248 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2249 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2250 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2251 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2252 VDD wake_up_sg a_10024_15996# VDD sg13g2_lv_pmos ad=0.2114p pd=1.54u as=0.2856p ps=2.36u w=0.84u l=0.13u
N2253 sg13g2_a21o_1_0.A2 sg13g2_buf_1_5.X VDD VDD sg13g2_lv_pmos ad=0.2128p pd=1.5u as=0.3808p ps=2.92u w=1.12u l=0.13u
N2254 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2255 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2256 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2257 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2258 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2259 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2260 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2261 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2262 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2263 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2264 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2265 a_12777_14531# a_12420_14488# VDD VDD sg13g2_lv_pmos ad=63f pd=0.72u as=0.1563p ps=1.22u w=0.42u l=0.13u
N2266 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2267 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2268 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2269 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2270 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2271 a_12134_14922# sg13g2_nor2b_1_0.Y VDD VDD sg13g2_lv_pmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
N2272 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2273 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2274 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2275 sg13g2_nor2_1_0.A a_10024_15996# VDD VDD sg13g2_lv_pmos ad=0.42p pd=2.99u as=0.2114p ps=1.54u w=1.12u l=0.13u
N2276 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2277 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2278 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2279 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2280 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2281 a_14314_15964# a_14757_16007# a_14697_16043# VDD sg13g2_lv_pmos ad=79.8f pd=0.8u as=63f ps=0.72u w=0.42u l=0.13u
N2282 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2283 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2284 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2285 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2286 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2287 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2288 sg13g2_a21o_1_1.A2 sg13g2_inv_2_1.A VDD VDD sg13g2_lv_pmos ad=0.2128p pd=1.5u as=0.3808p ps=2.92u w=1.12u l=0.13u
N2289 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2290 a_14061_12256# sg13g2_buf_1_4.A VDD VDD sg13g2_lv_pmos ad=0.1596p pd=1.22u as=0.2856p ps=2.36u w=0.84u l=0.13u
N2291 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2292 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2293 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2294 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2295 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2296 sg13g2_inv_2_1.A a_17800_15272# VSS VSS sg13g2_lv_nmos ad=0.2886p pd=2.26u as=0.14875p ps=1.16u w=0.74u l=0.13u
N2297 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2298 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2299 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2300 adc_start a_17128_13760# VSS VSS sg13g2_lv_nmos ad=0.2886p pd=2.26u as=0.14875p ps=1.16u w=0.74u l=0.13u
N2301 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2302 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2303 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2304 a_14949_13701# sg13g2_dfrbpq_1_0.CLK a_15409_13743# VSS sg13g2_lv_nmos ad=0.2516p pd=2.16u as=0.31732p ps=1.805u w=0.74u l=0.13u
N2305 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2306 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2307 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2308 a_14998_16742# sg13g2_a22oi_1_0.B2 VSS VSS sg13g2_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.15u
N2309 a_11076_16000# a_11050_15964# VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0.36237p ps=2.605u w=1u l=0.13u
N2310 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2311 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2312 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2313 a_11302_16421# sg13g2_inv_1_0.Y VSS VSS sg13g2_lv_nmos ad=37.8f pd=0.6u as=0.1701p ps=1.65u w=0.42u l=0.13u
N2314 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2315 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2316 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2317 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2318 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2319 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2320 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2321 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2322 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2323 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2324 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2325 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2326 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2327 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2328 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2329 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2330 sg13g2_a22oi_1_0.B2 a_15976_25068# VSS VSS sg13g2_lv_nmos ad=0.2886p pd=2.26u as=0.14875p ps=1.16u w=0.74u l=0.13u
N2331 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2332 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2333 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2334 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2335 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2336 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2337 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2338 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2339 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2340 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2341 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2342 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2343 VSS sg13g2_a21oi_1_0.A2 a_13601_16344# VSS sg13g2_lv_nmos ad=0.2516p pd=2.16u as=0.1406p ps=1.12u w=0.74u l=0.13u
N2344 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2345 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2346 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2347 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2348 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2349 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2350 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2351 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2352 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2353 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2354 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2355 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2356 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2357 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2358 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2359 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2360 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2361 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2362 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2363 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2364 a_11050_15964# a_11493_16007# a_10790_16434# VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0.1296p ps=1.52u w=0.42u l=0.13u
N2365 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2366 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2367 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2368 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2369 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2370 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2371 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2372 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2373 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2374 VSS sg13g2_a21oi_1_0.A2 a_14235_17564# VSS sg13g2_lv_nmos ad=0.14505p pd=1.15u as=0.187p ps=1.78u w=0.55u l=0.13u
N2375 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2376 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2377 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2378 sg13g2_nor2_1_0.B a_13002_15996# VDD VDD sg13g2_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
N2379 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2380 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2381 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2382 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2383 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2384 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2385 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2386 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2387 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2388 a_12326_16746# sg13g2_dfrbpq_1_6.D VDD VDD sg13g2_lv_pmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
N2389 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2390 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2391 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2392 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2393 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2394 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2395 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2396 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2397 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2398 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2399 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2400 a_13297_14837# a_12837_14495# a_12939_14495# VSS sg13g2_lv_nmos ad=0.31732p pd=1.805u as=0.2516p ps=2.16u w=0.74u l=0.13u
N2401 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2402 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2403 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2404 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2405 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2406 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2407 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2408 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2409 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2410 VDD uart_busy a_15976_25068# VDD sg13g2_lv_pmos ad=0.2114p pd=1.54u as=0.2856p ps=2.36u w=0.84u l=0.13u
N2411 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2412 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2413 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2414 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2415 sg13g2_a21oi_1_0.A2 a_13960_25068# VDD VDD sg13g2_lv_pmos ad=0.42p pd=2.99u as=0.2114p ps=1.54u w=1.12u l=0.13u
N2416 VSS sg13g2_inv_1_0.Y a_10884_16434# VSS sg13g2_lv_nmos ad=0.1626p pd=1.415u as=60.89999f ps=0.71u w=0.42u l=0.13u
N2417 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2418 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2419 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2420 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2421 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2422 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2423 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2424 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2425 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2426 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2427 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2428 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2429 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2430 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2431 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2432 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2433 a_11953_15998# a_11493_16007# a_11595_16007# VDD sg13g2_lv_pmos ad=0.41165p pd=2.12u as=0.3864p ps=2.93u w=1.12u l=0.13u
N2434 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2435 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2436 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2437 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2438 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2439 a_12335_16357# a_11493_16007# a_11076_16000# VDD sg13g2_lv_pmos ad=0.2048p pd=1.63u as=0.34p ps=2.68u w=1u l=0.13u
N2440 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2441 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2442 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2443 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2444 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2445 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2446 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2447 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2448 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2449 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2450 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2451 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2452 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2453 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2454 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2455 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2456 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2457 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2458 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2459 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2460 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2461 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2462 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2463 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2464 a_14757_16007# sg13g2_dfrbpq_1_0.CLK a_15217_15998# VDD sg13g2_lv_pmos ad=0.4088p pd=2.97u as=0.41165p ps=2.12u w=1.12u l=0.13u
N2465 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2466 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2467 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2468 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2469 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2470 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2471 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2472 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2473 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2474 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2475 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2476 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2477 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2478 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2479 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2480 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2481 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2482 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2483 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2484 a_12394_14452# a_12837_14495# a_12134_14922# VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0.1296p ps=1.52u w=0.42u l=0.13u
N2485 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2486 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2487 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2488 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2489 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2490 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2491 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2492 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2493 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2494 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2495 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2496 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2497 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2498 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2499 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2500 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2501 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2502 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2503 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2504 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2505 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2506 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2507 VSS a_13459_12404# sg13g2_a21o_1_0.X VSS sg13g2_lv_nmos ad=0.15745p pd=1.175u as=0.2351p ps=2.16u w=0.74u l=0.13u
N2508 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2509 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2510 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2511 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2512 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2513 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2514 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2515 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2516 a_13679_14845# a_12837_14495# a_12420_14488# VDD sg13g2_lv_pmos ad=0.2048p pd=1.63u as=0.34p ps=2.68u w=1u l=0.13u
N2517 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2518 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2519 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2520 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2521 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2522 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2523 VSS a_15791_13799# a_16458_14020# VSS sg13g2_lv_nmos ad=0.1406p pd=1.12u as=0.2516p ps=2.16u w=0.74u l=0.13u
N2524 VDD sg13g2_a21oi_1_0.A1 a_13499_15996# VDD sg13g2_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
N2525 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2526 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2527 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2528 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2529 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2530 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2531 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2532 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2533 VDD sg13g2_buf_1_5.X a_14061_12256# VDD sg13g2_lv_pmos ad=0.1918p pd=1.5u as=0.1596p ps=1.22u w=0.84u l=0.13u
N2534 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2535 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2536 a_12357_13701# sg13g2_dfrbpq_1_0.CLK a_12817_13743# VSS sg13g2_lv_nmos ad=0.2516p pd=2.16u as=0.31732p ps=1.805u w=0.74u l=0.13u
N2537 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2538 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2539 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2540 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2541 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2542 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2543 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2544 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2545 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2546 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2547 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2548 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2549 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2550 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2551 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2552 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2553 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2554 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2555 VSS sg13g2_buf_1_4.A a_13768_10736# VSS sg13g2_lv_nmos ad=0.14875p pd=1.16u as=0.187p ps=1.78u w=0.55u l=0.13u
N2556 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2557 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2558 tx_start a_14248_23556# VSS VSS sg13g2_lv_nmos ad=0.2886p pd=2.26u as=0.14875p ps=1.16u w=0.74u l=0.13u
N2559 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2560 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2561 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2562 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2563 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2564 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2565 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2566 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2567 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2568 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2569 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2570 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2571 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2572 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2573 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2574 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2575 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2576 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2577 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2578 VSS a_12335_16357# a_13002_15996# VSS sg13g2_lv_nmos ad=0.1406p pd=1.12u as=0.2516p ps=2.16u w=0.74u l=0.13u
N2579 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2580 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2581 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2582 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2583 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2584 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2585 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2586 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2587 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2588 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2589 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2590 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2591 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2592 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2593 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2594 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2595 a_14246_15234# sg13g2_dfrbpq_1_3.D VDD VDD sg13g2_lv_pmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
N2596 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2597 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2598 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2599 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2600 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2601 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2602 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2603 a_13029_16725# sg13g2_dfrbpq_1_0.CLK a_13489_16767# VSS sg13g2_lv_nmos ad=0.2516p pd=2.16u as=0.31732p ps=1.805u w=0.74u l=0.13u
N2604 a_15993_15549# a_15051_15356# a_15791_15311# VDD sg13g2_lv_pmos ad=93.45f pd=0.865u as=0.2048p ps=1.63u w=0.42u l=0.13u
N2605 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2606 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2607 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2608 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2609 a_10884_16434# sg13g2_dfrbpq_1_4.D a_10790_16434# VSS sg13g2_lv_nmos ad=60.89999f pd=0.71u as=0.1428p ps=1.52u w=0.42u l=0.13u
N2610 a_12228_13735# a_12459_13844# a_11914_13945# VSS sg13g2_lv_nmos ad=0.2373p pd=1.97u as=79.8f ps=0.8u w=0.42u l=0.13u
N2611 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2612 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2613 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2614 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2615 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2616 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2617 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2618 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2619 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2620 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2621 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2622 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2623 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2624 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2625 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2626 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2627 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2628 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2629 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2630 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2631 a_16735_16388# sg13g2_dfrbpq_1_5.Q VSS VSS sg13g2_lv_nmos ad=0.13875p pd=1.115u as=0.2553p ps=2.17u w=0.74u l=0.13u
N2632 VDD sg13g2_a21oi_1_0.A1 a_14248_23556# VDD sg13g2_lv_pmos ad=0.2114p pd=1.54u as=0.2856p ps=2.36u w=0.84u l=0.13u
N2633 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2634 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2635 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2636 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2637 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2638 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2639 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2640 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2641 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2642 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2643 VDD a_13871_16823# a_14128_16966# VDD sg13g2_lv_pmos ad=0.4659p pd=3.65u as=79.8f ps=0.8u w=0.42u l=0.13u
N2644 a_11914_13945# a_12357_13701# a_12297_14113# VDD sg13g2_lv_pmos ad=79.8f pd=0.8u as=63f ps=0.72u w=0.42u l=0.13u
N2645 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2646 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2647 VSS sg13g2_dfrbpq_1_1.Q a_17128_13760# VSS sg13g2_lv_nmos ad=0.14875p pd=1.16u as=0.187p ps=1.78u w=0.55u l=0.13u
N2648 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2649 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2650 a_14246_13722# a_15051_13844# a_14506_13945# VDD sg13g2_lv_pmos ad=0.1428p pd=1.52u as=79.8f ps=0.8u w=0.42u l=0.13u
N2651 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2652 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2653 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2654 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2655 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2656 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2657 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2658 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2659 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2660 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2661 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2662 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2663 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2664 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2665 a_16108_14037# a_16048_13942# a_15993_14037# VDD sg13g2_lv_pmos ad=0.204p pd=1.835u as=93.45f ps=0.865u w=0.42u l=0.13u
N2666 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2667 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2668 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2669 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2670 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2671 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2672 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2673 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2674 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2675 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2676 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2677 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2678 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2679 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2680 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2681 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2682 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2683 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2684 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2685 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2686 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2687 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2688 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2689 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2690 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2691 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2692 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2693 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2694 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2695 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2696 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2697 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2698 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2699 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2700 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2701 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2702 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2703 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2704 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2705 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2706 sg13g2_buf_1_0.A a_14346_14484# VDD VDD sg13g2_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
N2707 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2708 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2709 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2710 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2711 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2712 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2713 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2714 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2715 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2716 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2717 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2718 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2719 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2720 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2721 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2722 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2723 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2724 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2725 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2726 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2727 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2728 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2729 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2730 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2731 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2732 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2733 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2734 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2735 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2736 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2737 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2738 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2739 a_12586_16969# a_13029_16725# a_12969_17137# VDD sg13g2_lv_pmos ad=79.8f pd=0.8u as=63f ps=0.72u w=0.42u l=0.13u
N2740 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2741 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2742 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2743 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2744 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2745 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2746 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2747 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2748 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2749 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2750 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2751 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2752 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2753 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2754 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2755 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2756 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2757 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2758 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2759 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2760 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2761 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2762 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2763 a_12228_13735# a_11940_14040# a_12166_13735# VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=37.8f ps=0.6u w=0.42u l=0.13u
N2764 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2765 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2766 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2767 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2768 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2769 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2770 VSS a_13199_13799# a_13866_14020# VSS sg13g2_lv_nmos ad=0.1406p pd=1.12u as=0.2516p ps=2.16u w=0.74u l=0.13u
N2771 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2772 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2773 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2774 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2775 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2776 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2777 sg13g2_nor2_1_0.Y sg13g2_nor2_1_0.B a_12650_15532# VDD sg13g2_lv_pmos ad=0.3808p pd=2.92u as=0.1176p ps=1.33u w=1.12u l=0.13u
N2778 sg13g2_buf_1_0.A a_14346_14484# VSS VSS sg13g2_lv_nmos ad=0.2516p pd=2.16u as=0.1406p ps=1.12u w=0.74u l=0.13u
N2779 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2780 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2781 sg13g2_dfrbpq_1_6.D sg13g2_o21ai_1_0.B1 a_14998_16742# VSS sg13g2_lv_nmos ad=0.2516p pd=2.16u as=0.1406p ps=1.12u w=0.74u l=0.15u
N2782 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2783 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2784 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2785 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2786 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2787 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2788 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2789 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2790 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2791 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2792 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2793 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2794 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2795 a_12335_16357# a_11493_16007# a_12241_16357# VSS sg13g2_lv_nmos ad=0.12665p pd=1.145u as=0.1428p ps=1.52u w=0.42u l=0.13u
N2796 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2797 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2798 a_12592_16238# sg13g2_inv_1_0.Y a_12652_16119# VDD sg13g2_lv_pmos ad=79.8f pd=0.8u as=0.204p ps=1.835u w=0.42u l=0.13u
N2799 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2800 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2801 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2802 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2803 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2804 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2805 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2806 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2807 sg13g2_inv_1_1.Y sg13g2_inv_1_1.A VSS VSS sg13g2_lv_nmos ad=0.2516p pd=2.16u as=0.2516p ps=2.16u w=0.74u l=0.13u
N2808 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2809 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2810 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2811 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2812 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2813 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2814 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2815 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2816 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2817 a_12420_14488# a_12939_14495# a_13679_14845# VSS sg13g2_lv_nmos ad=0.3473p pd=2.71u as=0.12665p ps=1.145u w=0.74u l=0.13u
N2818 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2819 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2820 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2821 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2822 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2823 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2824 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2825 VSS sg13g2_inv_1_0.Y a_14340_15234# VSS sg13g2_lv_nmos ad=0.1626p pd=1.415u as=60.89999f ps=0.71u w=0.42u l=0.13u
N2826 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2827 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2828 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2829 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2830 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2831 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2832 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2833 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2834 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2835 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2836 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2837 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2838 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2839 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2840 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2841 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2842 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2843 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2844 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2845 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2846 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2847 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2848 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2849 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2850 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2851 VSS a_13871_16823# a_14538_17044# VSS sg13g2_lv_nmos ad=0.1406p pd=1.12u as=0.2516p ps=2.16u w=0.74u l=0.13u
N2852 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2853 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2854 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2855 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2856 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2857 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2858 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2859 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2860 a_13199_13799# a_12357_13701# a_11940_14040# VDD sg13g2_lv_pmos ad=0.2048p pd=1.63u as=0.34p ps=2.68u w=1u l=0.13u
N2861 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2862 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2863 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2864 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2865 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2866 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2867 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2868 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2869 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2870 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2871 VSS sg13g2_buf_1_0.A a_14440_5412# VSS sg13g2_lv_nmos ad=0.14875p pd=1.16u as=0.187p ps=1.78u w=0.55u l=0.13u
N2872 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2873 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2874 VSS sg13g2_o21ai_1_0.A1 a_14998_16742# VSS sg13g2_lv_nmos ad=0.1406p pd=1.12u as=0.2516p ps=2.16u w=0.74u l=0.15u
N2875 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2876 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2877 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2878 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2879 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2880 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2881 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2882 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2883 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2884 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2885 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2886 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2887 a_14506_13945# a_14949_13701# a_14889_14113# VDD sg13g2_lv_pmos ad=79.8f pd=0.8u as=63f ps=0.72u w=0.42u l=0.13u
N2888 a_16048_13942# a_15791_13799# a_16210_13722# VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=37.8f ps=0.6u w=0.42u l=0.13u
N2889 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2890 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2891 VSS clk a_7816_15996# VSS sg13g2_lv_nmos ad=0.14875p pd=1.16u as=0.187p ps=1.78u w=0.55u l=0.13u
N2892 VDD a_15599_16357# a_16266_15996# VDD sg13g2_lv_pmos ad=0.2128p pd=1.5u as=0.3864p ps=2.93u w=1.12u l=0.13u
N2893 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2894 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2895 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2896 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2897 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2898 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2899 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2900 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2901 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2902 a_13029_16725# sg13g2_dfrbpq_1_0.CLK a_13489_17042# VDD sg13g2_lv_pmos ad=0.4088p pd=2.97u as=0.41165p ps=2.12u w=1.12u l=0.13u
N2903 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2904 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2905 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2906 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2907 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2908 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2909 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2910 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2911 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2912 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2913 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2914 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2915 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2916 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2917 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2918 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2919 a_13516_14037# a_13456_13942# a_13401_14037# VDD sg13g2_lv_pmos ad=0.204p pd=1.835u as=93.45f ps=0.865u w=0.42u l=0.13u
N2920 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2921 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2922 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2923 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2924 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2925 a_14148_16434# sg13g2_inv_1_1.Y a_14054_16434# VSS sg13g2_lv_nmos ad=60.89999f pd=0.71u as=0.1428p ps=1.52u w=0.42u l=0.13u
N2926 a_16735_15972# sg13g2_a22oi_1_0.B2 sg13g2_inv_1_1.A VDD sg13g2_lv_pmos ad=0.2744p pd=1.61u as=0.2128p ps=1.5u w=1.12u l=0.13u
N2927 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2928 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2929 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2930 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2931 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2932 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2933 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2934 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2935 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2936 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2937 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2938 sg13g2_nor2_1_0.Y sg13g2_nor2_1_0.A VSS VSS sg13g2_lv_nmos ad=0.1406p pd=1.12u as=0.2516p ps=2.16u w=0.74u l=0.13u
N2939 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2940 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2941 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2942 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2943 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2944 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2945 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2946 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2947 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2948 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2949 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2950 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2951 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2952 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2953 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2954 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2955 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2956 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2957 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2958 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2959 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2960 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2961 a_12420_16746# sg13g2_dfrbpq_1_6.D a_12326_16746# VSS sg13g2_lv_nmos ad=60.89999f pd=0.71u as=0.1428p ps=1.52u w=0.42u l=0.13u
N2962 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2963 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2964 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2965 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2966 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2967 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2968 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2969 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2970 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2971 VDD a_15599_16357# a_15856_16238# VDD sg13g2_lv_pmos ad=0.4659p pd=3.65u as=79.8f ps=0.8u w=0.42u l=0.13u
N2972 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2973 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2974 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2975 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2976 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2977 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2978 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2979 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2980 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2981 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2982 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2983 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2984 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2985 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2986 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N2987 a_12326_16746# a_13131_16868# a_12586_16969# VDD sg13g2_lv_pmos ad=0.1428p pd=1.52u as=79.8f ps=0.8u w=0.42u l=0.13u
N2988 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2989 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2990 a_13702_12532# sg13g2_a21o_1_0.A2 VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0.19p ps=1.38u w=1u l=0.13u
N2991 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2992 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2993 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2994 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2995 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2996 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N2997 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N2998 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N2999 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3000 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3001 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3002 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3003 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3004 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3005 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3006 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3007 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3008 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3009 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3010 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3011 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3012 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3013 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3014 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3015 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3016 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3017 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3018 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3019 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3020 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3021 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3022 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3023 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3024 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3025 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3026 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3027 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3028 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3029 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3030 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3031 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3032 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3033 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3034 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3035 VDD a_12335_16357# a_12592_16238# VDD sg13g2_lv_pmos ad=0.4659p pd=3.65u as=79.8f ps=0.8u w=0.42u l=0.13u
N3036 VDD sg13g2_dfrbpq_1_3.Q a_16294_14484# VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0.2125p ps=1.425u w=1u l=0.13u
N3037 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3038 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3039 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3040 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3041 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3042 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3043 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3044 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3045 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3046 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3047 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3048 a_14098_14922# sg13g2_inv_1_0.Y VSS VSS sg13g2_lv_nmos ad=37.8f pd=0.6u as=79.8f ps=0.8u w=0.42u l=0.13u
N3049 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3050 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3051 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3052 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3053 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3054 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3055 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3056 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3057 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3058 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3059 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3060 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3061 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3062 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3063 VDD sg13g2_buf_1_5.X sg13g2_a21o_1_0.A2 VDD sg13g2_lv_pmos ad=0.3864p pd=2.93u as=0.2128p ps=1.5u w=1.12u l=0.13u
N3064 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3065 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3066 a_14566_16421# sg13g2_inv_1_0.Y VSS VSS sg13g2_lv_nmos ad=37.8f pd=0.6u as=0.1701p ps=1.65u w=0.42u l=0.13u
N3067 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3068 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3069 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3070 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3071 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3072 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3073 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3074 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3075 a_15791_13799# a_14949_13701# a_14532_14040# VDD sg13g2_lv_pmos ad=0.2048p pd=1.63u as=0.34p ps=2.68u w=1u l=0.13u
N3076 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3077 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3078 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3079 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3080 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3081 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3082 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3083 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3084 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3085 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3086 sg13g2_buf_1_6.X a_8968_13760# VSS VSS sg13g2_lv_nmos ad=0.2886p pd=2.26u as=0.14875p ps=1.16u w=0.74u l=0.13u
N3087 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3088 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3089 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3090 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3091 a_16048_15454# sg13g2_inv_1_0.Y a_16108_15549# VDD sg13g2_lv_pmos ad=79.8f pd=0.8u as=0.204p ps=1.835u w=0.42u l=0.13u
N3092 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3093 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3094 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3095 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3096 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3097 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3098 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3099 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3100 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3101 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3102 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3103 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3104 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3105 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3106 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3107 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3108 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3109 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3110 a_13456_13942# a_13199_13799# a_13618_13722# VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=37.8f ps=0.6u w=0.42u l=0.13u
N3111 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3112 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3113 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3114 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3115 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3116 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3117 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3118 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3119 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3120 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3121 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3122 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3123 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3124 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3125 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3126 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3127 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3128 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3129 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3130 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3131 sg13g2_inv_1_1.Y sg13g2_inv_1_1.A VDD VDD sg13g2_lv_pmos ad=0.3808p pd=2.92u as=0.3808p ps=2.92u w=1.12u l=0.13u
N3132 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3133 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3134 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3135 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3136 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3137 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3138 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3139 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3140 sg13g2_dfrbpq_1_3.Q a_16458_15532# VSS VSS sg13g2_lv_nmos ad=0.2516p pd=2.16u as=0.1406p ps=1.12u w=0.74u l=0.13u
N3141 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3142 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3143 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3144 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3145 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3146 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3147 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3148 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3149 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3150 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3151 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3152 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3153 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3154 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3155 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3156 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3157 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3158 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3159 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3160 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3161 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3162 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3163 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3164 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3165 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3166 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3167 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3168 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3169 a_15599_16357# a_14757_16007# a_14340_16000# VDD sg13g2_lv_pmos ad=0.2048p pd=1.63u as=0.34p ps=2.68u w=1u l=0.13u
N3170 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3171 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3172 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3173 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3174 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3175 a_12650_15532# sg13g2_nor2_1_0.A VDD VDD sg13g2_lv_pmos ad=0.1176p pd=1.33u as=0.4032p ps=2.96u w=1.12u l=0.13u
N3176 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3177 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3178 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3179 a_14128_16966# a_13871_16823# a_14290_16746# VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=37.8f ps=0.6u w=0.42u l=0.13u
N3180 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3181 sg13g2_dfrbpq_1_6.D sg13g2_a22oi_1_0.B2 a_15096_17064# VDD sg13g2_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.15u
N3182 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3183 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3184 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3185 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3186 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3187 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3188 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3189 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3190 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3191 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3192 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3193 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3194 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3195 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3196 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3197 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3198 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3199 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3200 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3201 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3202 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3203 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3204 a_13871_16823# a_13029_16725# a_12612_17064# VDD sg13g2_lv_pmos ad=0.2048p pd=1.63u as=0.34p ps=2.68u w=1u l=0.13u
N3205 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3206 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3207 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3208 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3209 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3210 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3211 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3212 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3213 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3214 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3215 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3216 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3217 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3218 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3219 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3220 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3221 a_13401_14037# a_12459_13844# a_13199_13799# VDD sg13g2_lv_pmos ad=93.45f pd=0.865u as=0.2048p ps=1.63u w=0.42u l=0.13u
N3222 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3223 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3224 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3225 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3226 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3227 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3228 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3229 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3230 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3231 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3232 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3233 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3234 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3235 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3236 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3237 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3238 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3239 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3240 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3241 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3242 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3243 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3244 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3245 a_16294_14484# sg13g2_a21o_1_1.A2 VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0.19p ps=1.38u w=1u l=0.13u
N3246 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3247 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3248 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3249 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3250 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3251 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3252 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3253 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3254 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3255 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3256 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3257 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3258 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3259 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3260 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3261 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3262 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3263 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3264 VSS sg13g2_inv_2_1.A sg13g2_a21o_1_1.A2 VSS sg13g2_lv_nmos ad=0.2516p pd=2.16u as=0.1406p ps=1.12u w=0.74u l=0.13u
N3265 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3266 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3267 VDD sg13g2_buf_1_4.A a_13768_10736# VDD sg13g2_lv_pmos ad=0.2114p pd=1.54u as=0.2856p ps=2.36u w=0.84u l=0.13u
N3268 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3269 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3270 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3271 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3272 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3273 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3274 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3275 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3276 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3277 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3278 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3279 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3280 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3281 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3282 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3283 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3284 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3285 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3286 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3287 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3288 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3289 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3290 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3291 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3292 a_13996_14607# a_13936_14726# a_13881_14607# VDD sg13g2_lv_pmos ad=0.204p pd=1.835u as=93.45f ps=0.865u w=0.42u l=0.13u
N3293 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3294 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3295 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3296 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3297 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3298 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3299 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3300 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3301 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3302 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3303 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3304 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3305 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3306 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3307 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3308 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3309 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3310 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3311 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3312 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3313 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3314 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3315 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3316 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3317 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3318 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3319 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3320 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3321 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3322 VDD adc_done a_17800_15272# VDD sg13g2_lv_pmos ad=0.2114p pd=1.54u as=0.2856p ps=2.36u w=0.84u l=0.13u
N3323 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3324 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3325 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3326 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3327 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3328 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3329 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3330 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3331 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3332 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3333 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3334 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3335 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3336 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3337 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3338 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3339 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3340 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3341 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3342 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3343 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3344 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3345 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3346 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3347 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3348 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3349 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3350 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3351 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3352 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3353 VDD sg13g2_inv_2_1.A a_16735_15972# VDD sg13g2_lv_pmos ad=0.3808p pd=2.92u as=0.2744p ps=1.61u w=1.12u l=0.13u
N3354 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3355 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3356 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3357 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3358 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3359 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3360 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3361 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3362 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3363 a_14340_15234# sg13g2_dfrbpq_1_3.D a_14246_15234# VSS sg13g2_lv_nmos ad=60.89999f pd=0.71u as=0.1428p ps=1.52u w=0.42u l=0.13u
N3364 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3365 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3366 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3367 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3368 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3369 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3370 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3371 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3372 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3373 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3374 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3375 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3376 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3377 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3378 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3379 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3380 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3381 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3382 VDD a_13459_12404# sg13g2_a21o_1_0.X VDD sg13g2_lv_pmos ad=0.3808p pd=2.92u as=0.3808p ps=2.92u w=1.12u l=0.13u
N3383 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3384 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3385 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3386 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3387 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3388 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3389 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3390 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3391 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3392 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3393 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3394 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3395 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3396 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3397 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3398 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3399 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3400 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3401 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3402 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3403 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3404 a_14437_17878# sg13g2_a21oi_1_0.A1 VSS VSS sg13g2_lv_nmos ad=0.1406p pd=1.12u as=0.14505p ps=1.15u w=0.74u l=0.13u
N3405 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3406 a_14246_13722# sg13g2_and2_1_0.X VDD VDD sg13g2_lv_pmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
N3407 VSS sg13g2_inv_1_0.Y a_14340_13722# VSS sg13g2_lv_nmos ad=0.1626p pd=1.415u as=60.89999f ps=0.71u w=0.42u l=0.13u
N3408 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3409 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3410 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3411 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3412 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3413 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3414 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3415 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3416 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3417 a_15993_14037# a_15051_13844# a_15791_13799# VDD sg13g2_lv_pmos ad=93.45f pd=0.865u as=0.2048p ps=1.63u w=0.42u l=0.13u
N3418 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3419 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3420 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3421 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3422 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3423 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3424 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3425 a_11364_16421# a_11076_16000# a_11302_16421# VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=37.8f ps=0.6u w=0.42u l=0.13u
N3426 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3427 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3428 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3429 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3430 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3431 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3432 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3433 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3434 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3435 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3436 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3437 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3438 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3439 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3440 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3441 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3442 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3443 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3444 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3445 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3446 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3447 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3448 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3449 a_13459_12404# sg13g2_buf_1_0.A VSS VSS sg13g2_lv_nmos ad=0.1216p pd=1.02u as=0.15745p ps=1.175u w=0.64u l=0.13u
N3450 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3451 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3452 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3453 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3454 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3455 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3456 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3457 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3458 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3459 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3460 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3461 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3462 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3463 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3464 a_12837_14495# sg13g2_dfrbpq_1_0.CLK a_13297_14837# VSS sg13g2_lv_nmos ad=0.2516p pd=2.16u as=0.31732p ps=1.805u w=0.74u l=0.13u
N3465 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3466 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3467 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3468 Timer_en a_13768_10736# VDD VDD sg13g2_lv_pmos ad=0.42p pd=2.99u as=0.2114p ps=1.54u w=1.12u l=0.13u
N3469 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3470 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3471 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3472 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3473 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3474 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3475 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3476 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3477 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3478 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3479 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3480 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3481 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3482 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3483 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3484 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3485 VDD sg13g2_inv_1_0.Y a_12134_14922# VDD sg13g2_lv_pmos ad=0.36237p pd=2.605u as=79.8f ps=0.8u w=0.42u l=0.13u
N3486 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3487 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3488 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3489 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3490 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3491 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3492 a_14054_16434# a_14859_16007# a_14314_15964# VDD sg13g2_lv_pmos ad=0.1428p pd=1.52u as=79.8f ps=0.8u w=0.42u l=0.13u
N3493 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3494 VDD sg13g2_inv_2_1.A sg13g2_a21o_1_1.A2 VDD sg13g2_lv_pmos ad=0.3864p pd=2.93u as=0.2128p ps=1.5u w=1.12u l=0.13u
N3495 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3496 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3497 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3498 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3499 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3500 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3501 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3502 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3503 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3504 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3505 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3506 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3507 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3508 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3509 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3510 sg13g2_buf_1_4.A a_13866_14020# VSS VSS sg13g2_lv_nmos ad=0.2516p pd=2.16u as=0.1406p ps=1.12u w=0.74u l=0.13u
N3511 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3512 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3513 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3514 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3515 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3516 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3517 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3518 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3519 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3520 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3521 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3522 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3523 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3524 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3525 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3526 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3527 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3528 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3529 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3530 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3531 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3532 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3533 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3534 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3535 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3536 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3537 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3538 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3539 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3540 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3541 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3542 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3543 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3544 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3545 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3546 VDD a_15791_15311# a_16458_15532# VDD sg13g2_lv_pmos ad=0.2128p pd=1.5u as=0.3864p ps=2.93u w=1.12u l=0.13u
N3547 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3548 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3549 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3550 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3551 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3552 a_11364_16421# a_11595_16007# a_11050_15964# VSS sg13g2_lv_nmos ad=0.2373p pd=1.97u as=79.8f ps=0.8u w=0.42u l=0.13u
N3553 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3554 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3555 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3556 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3557 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3558 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3559 a_10790_16434# sg13g2_dfrbpq_1_4.D VDD VDD sg13g2_lv_pmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
N3560 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3561 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3562 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3563 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3564 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3565 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3566 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3567 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3568 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3569 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3570 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3571 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3572 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3573 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3574 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3575 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3576 VDD sg13g2_inv_1_0.Y a_12326_16746# VDD sg13g2_lv_pmos ad=0.36237p pd=2.605u as=79.8f ps=0.8u w=0.42u l=0.13u
N3577 a_13881_14607# a_12939_14495# a_13679_14845# VDD sg13g2_lv_pmos ad=93.45f pd=0.865u as=0.2048p ps=1.63u w=0.42u l=0.13u
N3578 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3579 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3580 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3581 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3582 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3583 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3584 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3585 VDD sg13g2_o21ai_1_0.B1 sg13g2_dfrbpq_1_6.D VDD sg13g2_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.15u
N3586 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3587 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3588 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3589 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3590 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3591 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3592 a_14889_15625# a_14532_15552# VDD VDD sg13g2_lv_pmos ad=63f pd=0.72u as=0.1563p ps=1.22u w=0.42u l=0.13u
N3593 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3594 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3595 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3596 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3597 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3598 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3599 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3600 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3601 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3602 sc_en a_14440_5412# VDD VDD sg13g2_lv_pmos ad=0.42p pd=2.99u as=0.2114p ps=1.54u w=1.12u l=0.13u
N3603 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3604 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3605 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3606 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3607 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3608 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3609 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3610 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3611 VSS uart_busy a_15976_25068# VSS sg13g2_lv_nmos ad=0.14875p pd=1.16u as=0.187p ps=1.78u w=0.55u l=0.13u
N3612 a_11654_13722# sg13g2_a21o_1_0.X VDD VDD sg13g2_lv_pmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
N3613 sg13g2_a21oi_1_0.A2 a_13960_25068# VSS VSS sg13g2_lv_nmos ad=0.2886p pd=2.26u as=0.14875p ps=1.16u w=0.74u l=0.13u
N3614 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3615 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3616 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3617 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3618 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3619 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3620 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3621 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3622 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3623 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3624 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3625 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3626 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3627 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3628 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3629 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3630 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3631 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3632 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3633 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3634 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3635 VSS sg13g2_inv_1_0.Y a_14148_16434# VSS sg13g2_lv_nmos ad=0.1626p pd=1.415u as=60.89999f ps=0.71u w=0.42u l=0.13u
N3636 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3637 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3638 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3639 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3640 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3641 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3642 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3643 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3644 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3645 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3646 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3647 VSS wake_up_sg a_10024_15996# VSS sg13g2_lv_nmos ad=0.14875p pd=1.16u as=0.187p ps=1.78u w=0.55u l=0.13u
N3648 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3649 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3650 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3651 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3652 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3653 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3654 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3655 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3656 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3657 a_12708_14909# a_12939_14495# a_12394_14452# VSS sg13g2_lv_nmos ad=0.2373p pd=1.97u as=79.8f ps=0.8u w=0.42u l=0.13u
N3658 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3659 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3660 a_15096_17064# sg13g2_o21ai_1_0.A1 VDD VDD sg13g2_lv_pmos ad=0.2128p pd=1.5u as=0.3808p ps=2.92u w=1.12u l=0.15u
N3661 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3662 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3663 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3664 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3665 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3666 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3667 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3668 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3669 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3670 sg13g2_nor2_1_0.A a_10024_15996# VSS VSS sg13g2_lv_nmos ad=0.2886p pd=2.26u as=0.14875p ps=1.16u w=0.74u l=0.13u
N3671 VSS sg13g2_inv_1_0.Y a_12420_16746# VSS sg13g2_lv_nmos ad=0.1626p pd=1.415u as=60.89999f ps=0.71u w=0.42u l=0.13u
N3672 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3673 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3674 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3675 VDD uart_done a_13960_25068# VDD sg13g2_lv_pmos ad=0.2114p pd=1.54u as=0.2856p ps=2.36u w=0.84u l=0.13u
N3676 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3677 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3678 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3679 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3680 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3681 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3682 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3683 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3684 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3685 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3686 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3687 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3688 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3689 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3690 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3691 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3692 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3693 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3694 a_13499_15996# sg13g2_a21oi_1_0.A2 VDD VDD sg13g2_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
N3695 sg13g2_dfrbpq_1_1.Q a_16458_14020# VSS VSS sg13g2_lv_nmos ad=0.2516p pd=2.16u as=0.1406p ps=1.12u w=0.74u l=0.13u
N3696 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3697 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3698 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3699 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3700 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3701 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3702 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3703 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3704 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3705 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3706 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3707 VDD sg13g2_inv_1_0.Y a_11050_15964# VDD sg13g2_lv_pmos ad=0.1563p pd=1.22u as=0.147p ps=1.54u w=0.42u l=0.13u
N3708 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3709 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3710 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3711 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3712 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3713 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3714 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3715 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3716 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3717 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3718 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3719 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3720 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3721 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3722 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3723 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3724 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3725 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3726 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3727 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3728 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3729 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3730 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3731 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3732 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3733 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3734 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3735 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3736 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3737 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3738 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3739 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3740 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3741 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3742 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3743 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3744 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3745 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3746 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3747 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3748 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3749 sg13g2_nor2_1_0.B a_13002_15996# VSS VSS sg13g2_lv_nmos ad=0.2516p pd=2.16u as=0.1406p ps=1.12u w=0.74u l=0.13u
N3750 sg13g2_o21ai_1_0.B1 sg13g2_a21oi_1_0.A1 VDD VDD sg13g2_lv_pmos ad=0.2128p pd=1.5u as=0.2198p ps=1.53u w=1.12u l=0.13u
N3751 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3752 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3753 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3754 clk_gating_en a_14632_4688# VSS VSS sg13g2_lv_nmos ad=0.2886p pd=2.26u as=0.14875p ps=1.16u w=0.74u l=0.13u
N3755 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3756 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3757 VDD sg13g2_inv_1_0.Y a_10790_16434# VDD sg13g2_lv_pmos ad=0.36237p pd=2.605u as=79.8f ps=0.8u w=0.42u l=0.13u
N3758 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3759 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3760 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3761 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3762 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3763 VDD sg13g2_inv_1_0.Y a_14246_15234# VDD sg13g2_lv_pmos ad=0.36237p pd=2.605u as=79.8f ps=0.8u w=0.42u l=0.13u
N3764 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3765 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3766 VSS VDD VSS VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
N3767 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3768 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3769 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3770 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3771 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3772 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3773 sg13g2_dfrbpq_1_4.D sg13g2_nor2_1_0.Y VSS VSS sg13g2_lv_nmos ad=0.1406p pd=1.12u as=0.2516p ps=2.16u w=0.74u l=0.13u
N3774 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3775 VDD a_16051_14746# sg13g2_dfrbpq_1_3.D VDD sg13g2_lv_pmos ad=0.3808p pd=2.92u as=0.3808p ps=2.92u w=1.12u l=0.13u
N3776 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
N3777 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3778 VSS VDD VSS VSS sg13g2_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
N3779 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
N3780 VSS a_15856_16238# a_15505_16357# VSS sg13g2_lv_nmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
N3781 VDD VSS VDD VDD sg13g2_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
C0 a_17006_16388# sg13g2_dfrbpq_1_5.Q 0
C1 a_14235_17564# sg13g2_o21ai_1_0.B1 0.29113f
C2 a_13960_4782# a_14144_4782# 0.0524f
C3 a_14889_15625# sg13g2_inv_1_1.A 0
C4 a_17024_13854# VDD 0.06319f
C5 a_15791_13799# a_16051_14746# 0
C6 a_12459_13844# VDD 0.19509f
C7 a_12134_14922# a_12777_14531# 0.00801f
C8 a_12837_14495# a_13679_14845# 0.00307f
C9 a_12708_14909# a_12939_14495# 0.12701f
C10 uart_en sg13g2_buf_1_0.A 0.03977f
C11 a_13866_14020# sg13g2_inv_1_0.Y 0.01461f
C12 a_13002_15996# sg13g2_inv_1_1.Y 0
C13 adc_done sg13g2_a21o_1_1.A2 0
C14 sg13g2_dfrbpq_1_5.Q a_15680_16878# 0.01758f
C15 a_15051_15356# a_16048_15454# 0.02979f
C16 sg13g2_buf_1_0.A a_13576_4688# 0.2758f
C17 sg13g2_dfrbpq_1_6.D a_13864_16426# 0.00193f
C18 a_12612_17064# sg13g2_nor2_1_0.Y 0.00461f
C19 a_14340_16000# a_15599_16357# 0.01529f
C20 a_14757_16007# a_15856_16238# 0
C21 a_15993_14037# sg13g2_dfrbpq_1_1.Q 0
C22 a_13105_13799# a_12459_13844# 0.00647f
C23 a_13866_14020# a_13199_13799# 0.0894f
C24 uart_done a_13960_25068# 0.26647f
C25 a_12650_15532# sg13g2_nor2_1_0.Y 0.01296f
C26 a_13516_14037# VDD 0.00769f
C27 a_12900_16759# sg13g2_nor2_1_0.Y 0.0025f
C28 a_13679_14845# a_14346_14484# 0.0894f
C29 a_13936_14726# a_13585_14845# 0.008f
C30 sg13g2_buf_1_0.A a_13960_4572# 0.00147f
C31 a_13499_15996# sg13g2_a21oi_1_0.A2 0.07879f
C32 sg13g2_a22oi_1_0.B2 sg13g2_inv_1_1.Y 0.0025f
C33 a_15051_15356# a_15409_15255# 0.00104f
C34 a_14949_15213# a_15697_15311# 0.01058f
C35 a_16048_15454# a_16108_15549# 0.01042f
C36 a_15791_15311# a_16458_15532# 0.0894f
C37 sg13g2_inv_1_1.A a_12612_17064# 0
C38 a_14340_16000# sg13g2_dfrbpq_1_4.D 0
C39 a_16832_15366# sg13g2_inv_1_1.A 0.00394f
C40 sg13g2_nor2_1_0.A a_11493_16007# 0.00154f
C41 a_17024_13644# sg13g2_dfrbpq_1_1.Q 0.00102f
C42 sg13g2_a21oi_1_0.A1 a_13029_16725# 0.00184f
C43 a_13585_14845# sg13g2_buf_1_0.A 0
C44 a_12650_15532# sg13g2_inv_1_1.A 0
C45 a_15496_16668# sg13g2_dfrbpq_1_6.D 0.00618f
C46 a_9728_13854# VDD 0.10036f
C47 a_15051_15356# sg13g2_dfrbpq_1_0.CLK 0.04384f
C48 a_13960_25068# a_13856_25154# 0.00624f
C49 a_14506_15457# sg13g2_a21oi_1_0.A1 0
C50 adc_done a_25856_16668# 0
C51 a_15791_15311# a_16210_15234# 0.00174f
C52 a_16048_15454# a_15697_15311# 0.008f
C53 sg13g2_o21ai_1_0.A1 a_15496_16668# 0.00237f
C54 a_16266_15996# sg13g2_dfrbpq_1_3.Q 0.01003f
C55 a_14144_17938# sg13g2_a21oi_1_0.A2 0.00228f
C56 sg13g2_a22oi_1_0.B2 a_15916_16119# 0.00187f
C57 a_13401_14037# sg13g2_a21o_1_0.X 0
C58 a_14144_17594# VDD 0.08419f
C59 a_12326_16746# a_13871_16823# 0
C60 sg13g2_inv_1_1.A sg13g2_dfrbpq_1_5.Q 0.11359f
C61 sg13g2_a22oi_1_0.B2 a_15680_16668# 0
C62 sg13g2_nor2_1_0.A a_12136_16878# 0
C63 a_14073_17061# a_13871_16823# 0.00689f
C64 a_16108_15549# sg13g2_dfrbpq_1_0.CLK 0.00139f
C65 a_14061_12256# sg13g2_inv_1_0.Y 0
C66 a_12754_16434# sg13g2_nor2_1_0.Y 0
C67 adc_start a_17696_15156# 0
C68 a_13459_12404# a_13702_12532# 0.13617f
C69 sg13g2_dfrbpq_1_4.D sg13g2_a21oi_1_0.A2 0.00432f
C70 a_11848_15366# sg13g2_nor2_1_0.A 0.03085f
C71 a_13864_16082# a_14054_16434# 0.00201f
C72 a_14054_16434# a_13679_14845# 0
C73 sg13g2_a21oi_1_0.A1 a_11953_16349# 0
C74 a_12394_14452# VDD 0.10067f
C75 a_12326_16746# a_13489_17042# 0
C76 a_12612_17064# a_13131_16868# 0.34114f
C77 wake_up_sg VDD 1.55825f
C78 a_15697_15311# sg13g2_dfrbpq_1_0.CLK 0.00441f
C79 sg13g2_nor2b_1_0.Y sg13g2_nor2_1_0.Y 0.00972f
C80 a_13489_16767# a_12612_17064# 0.01835f
C81 a_12900_16759# a_13131_16868# 0.12701f
C82 a_13472_4572# VDD 0
C83 a_16430_14832# VDD 0
C84 sg13g2_dfrbpq_1_3.D a_16832_15366# 0
C85 a_14532_15552# sg13g2_o21ai_1_0.A1 0
C86 uart_busy tx_start 0.13424f
C87 a_13499_15996# VDD 0.26397f
C88 a_12900_16759# a_13489_16767# 0
C89 a_13936_14726# VDD 0.17826f
C90 sg13g2_dfrbpq_1_1.Q a_16832_15156# 0
C91 sg13g2_a22oi_1_0.B2 a_15505_16357# 0.00763f
C92 a_14949_15213# sg13g2_inv_2_1.A 0
C93 sg13g2_a22oi_1_0.B2 tx_start 0.05338f
C94 a_14949_15213# sg13g2_a22oi_1_0.B2 0.00126f
C95 a_14144_17938# VDD 0.00264f
C96 a_13192_12342# sg13g2_a21o_1_0.X 0.03677f
C97 a_15791_15311# sg13g2_o21ai_1_0.A1 0
C98 a_15599_16357# VDD 0.18329f
C99 sg13g2_dfrbpq_1_3.D a_14246_13722# 0.00156f
C100 sg13g2_dfrbpq_1_3.D sg13g2_dfrbpq_1_5.Q 0
C101 sg13g2_dfrbpq_1_0.CLK a_11493_16007# 0.27541f
C102 a_15217_15998# sg13g2_inv_1_0.Y 0.01659f
C103 sg13g2_buf_1_0.A VDD 2.76775f
C104 sg13g2_dfrbpq_1_6.D a_13871_16823# 0.02117f
C105 a_16048_15454# sg13g2_inv_2_1.A 0.00118f
C106 sg13g2_dfrbpq_1_1.Q a_16294_14484# 0.08523f
C107 sg13g2_o21ai_1_0.A1 a_13871_16823# 0
C108 a_14538_17044# a_14128_16966# 0.10373f
C109 a_14889_14113# sg13g2_dfrbpq_1_0.CLK 0
C110 a_16048_15454# sg13g2_a22oi_1_0.B2 0
C111 a_13105_13799# sg13g2_buf_1_0.A 0.00141f
C112 a_14889_15625# sg13g2_inv_1_0.Y 0
C113 a_13864_16082# sg13g2_inv_1_1.Y 0.04058f
C114 a_14061_12256# timer_done 0
C115 a_12326_16746# sg13g2_nor2_1_0.B 0
C116 sg13g2_dfrbpq_1_4.D VDD 0.42835f
C117 sg13g2_nor2_1_0.A a_11914_13945# 0
C118 a_14246_13722# a_14949_13701# 0.02454f
C119 sg13g2_dfrbpq_1_0.CLK a_13002_15996# 0.01183f
C120 a_11076_16000# a_11493_16007# 0.37384f
C121 sg13g2_inv_1_1.Y a_13679_14845# 0
C122 sg13g2_dfrbpq_1_6.D a_13489_17042# 0.00234f
C123 a_12136_16878# sg13g2_dfrbpq_1_0.CLK 0.00266f
C124 a_14340_16000# a_15680_16878# 0
C125 a_14757_16007# a_15496_16878# 0.00238f
C126 a_17128_13760# sg13g2_dfrbpq_1_0.CLK 0
C127 a_13777_16823# sg13g2_dfrbpq_1_6.D 0.00577f
C128 a_14538_17044# sg13g2_dfrbpq_1_0.CLK 0
C129 a_13601_16344# sg13g2_a21oi_1_0.A2 0.00205f
C130 a_14532_14040# a_15791_13799# 0.01529f
C131 sg13g2_dfrbpq_1_3.Q sg13g2_dfrbpq_1_1.Q 0.15484f
C132 sg13g2_buf_1_5.X Timer_en 0.02836f
C133 a_11848_15366# sg13g2_dfrbpq_1_0.CLK 0
C134 a_11364_16421# a_11595_16007# 0.12701f
C135 a_11493_16007# a_12335_16357# 0.00307f
C136 sg13g2_dfrbpq_1_3.D a_14820_13735# 0
C137 a_10790_16434# a_11433_16043# 0.00801f
C138 a_14538_17044# a_14290_16746# 0
C139 sg13g2_inv_2_1.A sg13g2_dfrbpq_1_0.CLK 0.0041f
C140 a_12136_16878# a_11076_16000# 0
C141 sg13g2_a22oi_1_0.B2 sg13g2_dfrbpq_1_0.CLK 0.22482f
C142 sg13g2_inv_1_0.Y a_12612_17064# 0.40714f
C143 a_12586_16969# a_13029_16725# 0.02242f
C144 sg13g2_dfrbpq_1_0.CLK a_12817_14018# 0.00251f
C145 sg13g2_nor2_1_0.A a_12420_14488# 0
C146 a_12046_15276# a_11493_16007# 0.00159f
C147 a_11848_15366# a_11076_16000# 0
C148 a_12900_16759# sg13g2_inv_1_0.Y 0.00396f
C149 a_15051_13844# a_15993_14037# 0
C150 a_14532_14040# a_14758_13735# 0.0052f
C151 a_14949_13701# a_14820_13735# 0.01562f
C152 a_12335_16357# a_13002_15996# 0.0894f
C153 a_12592_16238# a_12241_16357# 0.008f
C154 a_12650_15532# sg13g2_inv_1_0.Y 0.00356f
C155 timer_done sc_en 0.27424f
C156 sg13g2_dfrbpq_1_3.Q a_15801_16119# 0
C157 sg13g2_dfrbpq_1_6.D a_12592_16238# 0.0019f
C158 sc_en a_14632_4688# 0.04835f
C159 sg13g2_inv_1_1.A a_17696_15366# 0
C160 a_12228_13735# VDD 0.00693f
C161 sg13g2_nor2b_1_0.Y a_11595_16007# 0.00132f
C162 a_13864_16426# a_14054_16434# 0.00404f
C163 sg13g2_dfrbpq_1_5.Q sg13g2_inv_1_0.Y 0.00147f
C164 a_12241_16357# sg13g2_nor2_1_0.B 0
C165 a_16458_14020# a_17128_13760# 0
C166 a_14246_13722# sg13g2_inv_1_0.Y 0.11428f
C167 sg13g2_a21o_1_0.A2 sg13g2_buf_1_5.X 0.29471f
C168 a_12046_15276# a_12136_16878# 0
C169 sg13g2_and2_1_0.X a_14949_13701# 0.00142f
C170 a_14506_13945# a_15051_13844# 0.01f
C171 a_14340_16000# sg13g2_inv_1_1.A 0.00147f
C172 sg13g2_dfrbpq_1_6.D sg13g2_nor2_1_0.B 0.00235f
C173 sg13g2_inv_1_0.Y a_11364_16421# 0
C174 a_12046_15276# a_11848_15366# 0.01393f
C175 sg13g2_a21oi_1_0.A1 a_14757_16007# 0.00668f
C176 sg13g2_o21ai_1_0.B1 a_13871_16823# 0.00207f
C177 a_13480_10830# sg13g2_buf_1_0.A 0.00926f
C178 a_14340_13722# sg13g2_inv_1_0.Y 0
C179 a_15784_14570# VDD 0.16488f
C180 a_14820_13735# a_15409_13743# 0
C181 sg13g2_and2_1_0.X a_16048_13942# 0
C182 a_17024_13854# a_17128_13760# 0.00624f
C183 a_13601_16344# VDD 0
C184 a_13618_13722# a_13456_13942# 0.00188f
C185 a_15599_16357# a_16018_16434# 0.00174f
C186 a_14859_16007# a_15217_15998# 0.02138f
C187 a_13881_14607# VDD 0.00138f
C188 sg13g2_inv_1_0.Y a_12754_16434# 0.00114f
C189 sg13g2_a21oi_1_0.A1 a_15217_16349# 0
C190 sg13g2_a21oi_1_0.A1 a_14144_23642# 0.02298f
C191 a_15791_15311# a_16294_14484# 0
C192 sg13g2_nor2b_1_0.Y a_11940_14040# 0
C193 a_14152_5498# sg13g2_buf_1_0.A 0.01194f
C194 tx_start a_13960_25068# 0.00332f
C195 a_14532_15552# sg13g2_dfrbpq_1_3.Q 0
C196 a_15051_15356# a_15599_16357# 0
C197 a_14820_13735# sg13g2_inv_1_0.Y 0.00158f
C198 sg13g2_nor2b_1_0.Y sg13g2_inv_1_0.Y 0.18535f
C199 a_17006_16388# VDD 0
C200 sg13g2_and2_1_0.X a_15409_13743# 0
C201 sg13g2_buf_1_5.X sg13g2_a21o_1_0.X 0
C202 a_14061_12256# a_13866_14020# 0
C203 a_12459_13844# a_12817_14018# 0.02138f
C204 a_11654_13722# a_11748_13722# 0.00716f
C205 a_13702_12532# VDD 0.34097f
C206 a_15680_16878# VDD 0.07064f
C207 sg13g2_dfrbpq_1_0.CLK a_12420_14488# 0.10683f
C208 a_16840_13854# sg13g2_dfrbpq_1_0.CLK 0
C209 sg13g2_a21o_1_1.A2 a_16051_14746# 0.00145f
C210 a_15791_15311# sg13g2_dfrbpq_1_3.Q 0.00902f
C211 sg13g2_and2_1_0.X sg13g2_inv_1_0.Y 0.17346f
C212 sg13g2_dfrbpq_1_3.D a_14340_16000# 0
C213 a_13459_12404# sg13g2_inv_1_0.Y 0.00131f
C214 sg13g2_inv_1_0.Y a_11464_13644# 0.00247f
C215 sg13g2_inv_1_1.Y a_13996_14607# 0
C216 a_13459_12404# a_13199_13799# 0
C217 a_13864_16082# sg13g2_dfrbpq_1_0.CLK 0.01121f
C218 a_25856_11546# VDD 0.0583f
C219 sg13g2_dfrbpq_1_0.CLK a_13679_14845# 0.0105f
C220 a_10024_15996# VDD 0.26883f
C221 wake_up_sg a_11493_16007# 0
C222 sg13g2_nor2_1_0.Y VDD 0.44431f
C223 sg13g2_a21oi_1_0.A1 a_14314_15964# 0.00473f
C224 a_13131_16868# sg13g2_a21oi_1_0.A2 0.03088f
C225 a_11914_13945# a_12459_13844# 0.01f
C226 sg13g2_a21o_1_0.X a_11654_13722# 0.27608f
C227 a_14152_5842# VDD 0.00916f
C228 a_16266_15996# sg13g2_dfrbpq_1_0.CLK 0.00152f
C229 Timer_en a_14248_4688# 0.00655f
C230 a_12592_16238# a_12837_14495# 0
C231 a_12335_16357# a_12420_14488# 0
C232 reset VDD 1.34688f
C233 a_14859_16007# sg13g2_dfrbpq_1_5.Q 0
C234 a_14246_15234# VDD 0.79999f
C235 a_14336_5498# VDD 0.06961f
C236 a_16840_13854# a_16458_14020# 0.01012f
C237 a_13871_16823# a_14054_16434# 0
C238 sg13g2_nor2b_1_0.Y a_12134_14922# 0.27178f
C239 sg13g2_inv_1_0.Y a_11464_13854# 0.01456f
C240 sg13g2_inv_1_1.A VDD 0.53573f
C241 sg13g2_a21o_1_0.A2 sg13g2_a21o_1_0.X 0
C242 sg13g2_a21o_1_0.X a_11748_13722# 0
C243 sg13g2_nor2_1_0.B a_12837_14495# 0.0021f
C244 Timer_en a_14144_4572# 0.00131f
C245 a_14340_15234# VDD 0
C246 a_12459_13844# a_12420_14488# 0
C247 a_12357_13701# a_12837_14495# 0.00173f
C248 a_16840_13854# a_17024_13854# 0.0524f
C249 a_12420_16746# VDD 0
C250 sg13g2_dfrbpq_1_4.D a_11493_16007# 0.0131f
C251 a_16735_16388# sg13g2_a21o_1_1.A2 0
C252 a_15051_15356# a_15784_14570# 0
C253 a_14820_15247# VDD 0.00858f
C254 a_14340_16000# sg13g2_inv_1_0.Y 0.38254f
C255 a_14532_15552# sg13g2_inv_1_1.Y 0
C256 a_14506_15457# a_14314_15964# 0
C257 a_15856_16238# sg13g2_o21ai_1_0.A1 0
C258 sg13g2_inv_1_0.Y a_12646_14909# 0
C259 a_13456_13942# a_12837_14495# 0
C260 sg13g2_dfrbpq_1_4.D a_13002_15996# 0.01012f
C261 a_13131_16868# VDD 0.19128f
C262 a_12136_16878# sg13g2_dfrbpq_1_4.D 0
C263 sg13g2_a22oi_1_0.B2 a_15599_16357# 0.02317f
C264 a_16048_15454# sg13g2_dfrbpq_1_1.Q 0.00107f
C265 a_14628_16421# sg13g2_inv_1_0.Y 0.00138f
C266 sg13g2_dfrbpq_1_3.D VDD 0.48775f
C267 a_13489_16767# VDD 0
C268 a_13768_10736# a_14152_10736# 0.0015f
C269 sg13g2_a21oi_1_0.A1 a_14998_16742# 0.02723f
C270 sg13g2_inv_1_0.Y a_13585_14845# 0.00211f
C271 a_11848_15366# sg13g2_dfrbpq_1_4.D 0.0021f
C272 clk sg13g2_dfrbpq_1_0.CLK 0.06214f
C273 sg13g2_inv_1_1.A a_16735_15972# 0.1784f
C274 a_13199_13799# a_13585_14845# 0
C275 a_10884_16434# VDD 0
C276 a_13871_16823# sg13g2_inv_1_1.Y 0.001f
C277 a_13866_14020# a_14246_13722# 0
C278 sg13g2_inv_1_0.Y sg13g2_a21oi_1_0.A2 0.02943f
C279 a_15697_15311# a_15784_14570# 0
C280 a_14949_13701# VDD 0.2642f
C281 Timer_en adc_en 1.57613f
C282 a_11595_16007# VDD 0.18782f
C283 timer_done uart_en 0.76759f
C284 sg13g2_dfrbpq_1_0.CLK sg13g2_dfrbpq_1_1.Q 0.03476f
C285 sg13g2_buf_1_5.X sg13g2_buf_1_4.A 0.45745f
C286 timer_done a_13576_4688# 0
C287 uart_en a_14632_4688# 0.08855f
C288 a_16048_13942# VDD 0.16276f
C289 a_13777_16823# sg13g2_inv_1_1.Y 0.00102f
C290 sg13g2_dfrbpq_1_0.CLK a_13996_14607# 0.00143f
C291 a_14336_5842# a_14440_5412# 0
C292 sg13g2_dfrbpq_1_5.Q a_15784_14914# 0
C293 a_12394_14452# a_12420_14488# 0.36952f
C294 a_16210_13722# a_15697_13799# 0
C295 a_11953_15998# VDD 0.00645f
C296 a_11914_13945# sg13g2_buf_1_0.A 0
C297 a_15801_16119# sg13g2_dfrbpq_1_0.CLK 0.00134f
C298 Timer_en sg13g2_buf_1_4.A 0.00486f
C299 a_14152_5498# a_14336_5498# 0.0524f
C300 a_14532_15552# a_14949_15213# 0.3749f
C301 a_14246_15234# a_15051_15356# 0.097f
C302 timer_done a_13960_4572# 0
C303 a_15409_13743# VDD 0.00143f
C304 a_15051_15356# sg13g2_inv_1_1.A 0.02272f
C305 a_14248_4688# a_14144_4572# 0
C306 a_14235_17564# a_14144_17594# 0.00761f
C307 a_13192_12132# sg13g2_dfrbpq_1_0.CLK 0
C308 a_12837_14495# a_12939_14495# 0.47795f
C309 a_12420_14488# a_13936_14726# 0.00139f
C310 a_15496_16668# sg13g2_dfrbpq_1_0.CLK 0.00118f
C311 a_11940_14040# VDD 0.08626f
C312 a_15688_25154# VDD 0.1353f
C313 a_17024_13644# adc_start 0
C314 a_15791_13799# sg13g2_a21o_1_1.A2 0.00194f
C315 a_14246_15234# a_16108_15549# 0
C316 a_14532_15552# a_16048_15454# 0.00242f
C317 a_14949_15213# a_15791_15311# 0.00332f
C318 a_13105_13799# a_11940_14040# 0.43239f
C319 a_12817_13743# a_12357_13701# 0.02396f
C320 sg13g2_inv_1_0.Y VDD 10.0839f
C321 a_13866_14020# sg13g2_and2_1_0.X 0.01133f
C322 a_14340_16000# a_14859_16007# 0.34102f
C323 a_14757_16007# a_15217_16349# 0.02396f
C324 a_13499_15996# a_13864_16082# 0.01004f
C325 a_16458_14020# sg13g2_dfrbpq_1_1.Q 0.12431f
C326 a_9920_16082# sg13g2_dfrbpq_1_0.CLK 0.00209f
C327 a_16108_15549# sg13g2_inv_1_1.A 0.0031f
C328 a_13864_16082# a_13936_14726# 0
C329 a_13199_13799# VDD 0.18663f
C330 a_12420_14488# sg13g2_buf_1_0.A 0
C331 a_12837_14495# a_13297_14486# 0.01483f
C332 a_13936_14726# a_13679_14845# 0.34468f
C333 sg13g2_nor2_1_0.B sg13g2_inv_1_1.Y 0
C334 a_13105_13799# sg13g2_inv_1_0.Y 0.00532f
C335 sg13g2_a22oi_1_0.B2 a_15784_14570# 0
C336 sg13g2_buf_1_0.A a_13960_4782# 0.01025f
C337 sg13g2_a21o_1_0.A2 sg13g2_buf_1_4.A 0.5612f
C338 a_15791_15311# a_16048_15454# 0.34468f
C339 a_14532_15552# a_15409_15255# 0.01835f
C340 a_15051_15356# a_14820_15247# 0.12701f
C341 a_14628_16421# a_14859_16007# 0.12701f
C342 a_13105_13799# a_13199_13799# 0.28931f
C343 a_17024_13854# sg13g2_dfrbpq_1_1.Q 0.02574f
C344 sg13g2_dfrbpq_1_4.D a_12420_14488# 0
C345 a_15697_15311# sg13g2_inv_1_1.A 0
C346 sg13g2_nor2_1_0.A a_11050_15964# 0
C347 sg13g2_dfrbpq_1_3.D a_16018_16434# 0
C348 a_13679_14845# sg13g2_buf_1_0.A 0.00209f
C349 a_15496_16878# sg13g2_dfrbpq_1_6.D 0.02067f
C350 sg13g2_a21oi_1_0.A1 a_14073_17061# 0
C351 a_14532_15552# sg13g2_dfrbpq_1_0.CLK 0.09602f
C352 a_8776_13854# VDD 0.14617f
C353 a_11493_16007# sg13g2_nor2_1_0.Y 0
C354 a_14859_16007# sg13g2_a21oi_1_0.A2 0
C355 sg13g2_o21ai_1_0.A1 a_15496_16878# 0.00903f
C356 sg13g2_inv_2_1.A a_17006_16388# 0.00108f
C357 a_15856_16238# sg13g2_dfrbpq_1_3.Q 0.00142f
C358 a_15599_16357# a_16266_15996# 0.0894f
C359 sg13g2_dfrbpq_1_3.D a_15051_15356# 0.01234f
C360 a_13871_16823# a_14128_16966# 0.34468f
C361 a_13864_16082# sg13g2_dfrbpq_1_4.D 0.00113f
C362 a_12326_16746# a_12136_16668# 0.00404f
C363 a_14144_17938# a_14235_17564# 0
C364 a_12228_13735# a_11914_13945# 0.00463f
C365 sg13g2_nor2_1_0.A a_12592_16238# 0.00154f
C366 sg13g2_a21oi_1_0.A1 a_15096_17064# 0.00199f
C367 a_15791_15311# sg13g2_dfrbpq_1_0.CLK 0.00684f
C368 sg13g2_a22oi_1_0.B2 a_15680_16878# 0
C369 a_13459_12404# a_14061_12256# 0.00483f
C370 a_13002_15996# sg13g2_nor2_1_0.Y 0.05764f
C371 a_14061_12256# sg13g2_and2_1_0.X 0.10477f
C372 a_14757_16007# a_14314_15964# 0.02242f
C373 a_14949_15213# a_15051_13844# 0
C374 adc_en a_14248_4688# 0.02572f
C375 sg13g2_buf_1_4.A sg13g2_a21o_1_0.X 0
C376 sg13g2_dfrbpq_1_0.CLK a_13871_16823# 0
C377 sg13g2_nor2_1_0.A sg13g2_nor2_1_0.B 0.30504f
C378 a_12134_14922# VDD 0.79005f
C379 a_12326_16746# a_13029_16725# 0.02454f
C380 timer_done VDD 1.80756f
C381 a_14758_15247# sg13g2_dfrbpq_1_0.CLK 0
C382 a_14290_16746# a_13871_16823# 0.00174f
C383 a_13777_16823# a_14128_16966# 0.008f
C384 a_12900_16759# a_12612_17064# 0.43707f
C385 a_14632_4688# VDD 0.22656f
C386 sg13g2_nor2_1_0.A a_12357_13701# 0
C387 sg13g2_dfrbpq_1_3.D a_15697_15311# 0.02337f
C388 clk wake_up_sg 0.66497f
C389 sg13g2_a21oi_1_0.A1 a_12241_16357# 0
C390 a_12537_16119# VDD 0
C391 adc_en a_14144_4572# 0
C392 a_13489_17042# sg13g2_dfrbpq_1_0.CLK 0.00171f
C393 sg13g2_a21oi_1_0.A1 sg13g2_dfrbpq_1_6.D 0.15291f
C394 a_13297_14837# VDD 0.00223f
C395 a_14246_15234# sg13g2_a22oi_1_0.B2 0
C396 sg13g2_buf_1_6.X VDD 0.42191f
C397 a_25768_4782# VDD 0.13597f
C398 sg13g2_a21oi_1_0.A1 sg13g2_o21ai_1_0.A1 0.05349f
C399 sg13g2_a21o_1_1.A2 a_17696_15156# 0
C400 a_15791_15311# a_16458_14020# 0
C401 a_16458_15532# a_15791_13799# 0
C402 a_15697_15311# a_14949_13701# 0
C403 sg13g2_inv_2_1.A sg13g2_inv_1_1.A 0.69879f
C404 a_16832_15366# sg13g2_dfrbpq_1_5.Q 0.00116f
C405 a_14859_16007# VDD 0.19257f
C406 a_13777_16823# a_14290_16746# 0
C407 a_12777_14531# VDD 0
C408 a_25768_23986# VDD 0.00121f
C409 sg13g2_a22oi_1_0.B2 sg13g2_inv_1_1.A 0.27599f
C410 sg13g2_dfrbpq_1_0.CLK a_11050_15964# 0.0126f
C411 tx_start a_15872_25154# 0
C412 sg13g2_dfrbpq_1_6.D a_12136_16668# 0.00154f
C413 sg13g2_dfrbpq_1_1.Q a_16430_14832# 0
C414 a_15051_13844# sg13g2_dfrbpq_1_0.CLK 0.03561f
C415 a_15496_16878# sg13g2_o21ai_1_0.B1 0.01551f
C416 a_14188_17061# a_13871_16823# 0.00247f
C417 a_15697_15311# a_16048_13942# 0
C418 a_15051_15356# sg13g2_inv_1_0.Y 0.4257f
C419 a_11050_15964# a_11076_16000# 0.36952f
C420 a_16294_14484# a_16051_14746# 0.13617f
C421 sg13g2_dfrbpq_1_3.D a_14889_14113# 0
C422 sg13g2_dfrbpq_1_0.CLK a_12592_16238# 0.0107f
C423 sg13g2_dfrbpq_1_6.D a_13029_16725# 0.01883f
C424 a_13679_14845# a_13881_14607# 0.00689f
C425 a_13936_14726# a_13996_14607# 0.01042f
C426 a_16108_14037# sg13g2_dfrbpq_1_0.CLK 0.00139f
C427 a_14757_16007# a_14998_16742# 0.00108f
C428 a_12838_16759# sg13g2_dfrbpq_1_6.D 0
C429 sg13g2_o21ai_1_0.A1 a_13029_16725# 0
C430 a_14820_15247# sg13g2_a22oi_1_0.B2 0
C431 a_16108_15549# sg13g2_inv_1_0.Y 0.01227f
C432 a_15599_16357# sg13g2_dfrbpq_1_1.Q 0
C433 a_15051_13844# a_15409_14018# 0.02138f
C434 a_14246_13722# a_14340_13722# 0.00716f
C435 a_11076_16000# a_12592_16238# 0.00139f
C436 a_11493_16007# a_11595_16007# 0.47795f
C437 a_14506_15457# sg13g2_o21ai_1_0.A1 0
C438 sg13g2_dfrbpq_1_0.CLK sg13g2_nor2_1_0.B 0.13788f
C439 sg13g2_nor2b_1_0.Y a_12650_15532# 0
C440 sg13g2_dfrbpq_1_3.Q a_16051_14746# 0.01675f
C441 sg13g2_buf_1_0.A a_13996_14607# 0.00194f
C442 a_12586_16969# a_12326_16746# 0.75507f
C443 sg13g2_nor2_1_0.A a_12228_14922# 0
C444 sg13g2_dfrbpq_1_3.D sg13g2_inv_2_1.A 0.00235f
C445 a_15697_15311# sg13g2_inv_1_0.Y 0
C446 sg13g2_dfrbpq_1_3.D sg13g2_a22oi_1_0.B2 0
C447 sg13g2_dfrbpq_1_0.CLK a_12357_13701# 0.27179f
C448 sc_en uart_en 1.13309f
C449 a_15599_16357# a_15801_16119# 0.00689f
C450 a_15856_16238# a_15916_16119# 0.01042f
C451 a_12592_16238# a_12335_16357# 0.34468f
C452 wake_up_sg a_9920_16082# 0.02391f
C453 a_11493_16007# a_11953_15998# 0.01483f
C454 a_11076_16000# sg13g2_nor2_1_0.B 0
C455 a_14246_13722# a_14820_13735# 0.31978f
C456 a_16210_13722# adc_start 0
C457 a_12136_16878# a_11595_16007# 0
C458 sg13g2_nor2_1_0.Y a_12420_14488# 0
C459 sg13g2_a21oi_1_0.A1 sg13g2_o21ai_1_0.B1 0.15249f
C460 a_13866_14020# VDD 0.38905f
C461 a_13192_12132# sg13g2_buf_1_0.A 0.00234f
C462 a_11848_15366# a_11595_16007# 0
C463 a_15791_13799# a_15993_14037# 0.00689f
C464 a_14152_5498# timer_done 0.00315f
C465 sg13g2_dfrbpq_1_0.CLK a_13456_13942# 0.01698f
C466 a_12335_16357# sg13g2_nor2_1_0.B 0.0028f
C467 a_14506_13945# a_14532_14040# 0.36952f
C468 sg13g2_and2_1_0.X a_14246_13722# 0.27646f
C469 a_14340_16000# a_15217_15998# 0
C470 a_12228_13735# a_12166_13735# 0
C471 sg13g2_inv_1_0.Y a_11493_16007# 0.04385f
C472 sg13g2_a21oi_1_0.A1 a_12837_14495# 0
C473 a_13768_10736# sg13g2_buf_1_0.A 0.04455f
C474 a_12046_15276# sg13g2_nor2_1_0.B 0.06176f
C475 a_14889_14113# sg13g2_inv_1_0.Y 0
C476 a_14246_15234# a_13679_14845# 0
C477 a_17800_15272# a_17696_15366# 0.00624f
C478 sg13g2_and2_1_0.X a_14340_13722# 0
C479 a_15856_16238# a_15505_16357# 0.008f
C480 a_15784_14914# VDD 0.00332f
C481 sg13g2_inv_1_0.Y a_13002_15996# 0.0033f
C482 sg13g2_inv_1_1.A a_13679_14845# 0.0016f
C483 sg13g2_a21oi_1_0.A1 a_14566_16421# 0
C484 uart_busy a_15688_25154# 0.00537f
C485 a_9920_16082# sg13g2_dfrbpq_1_4.D 0
C486 a_14336_5842# sg13g2_buf_1_0.A 0
C487 sg13g2_inv_1_0.Y a_12136_16878# 0.00135f
C488 a_12586_16969# sg13g2_dfrbpq_1_6.D 0.01319f
C489 sg13g2_nor2_1_0.B a_12459_13844# 0.00155f
C490 a_15051_15356# a_14859_16007# 0
C491 a_15688_25498# a_15976_25068# 0
C492 sg13g2_and2_1_0.X a_14820_13735# 0.00326f
C493 a_14532_15552# sg13g2_buf_1_0.A 0
C494 a_11848_15366# sg13g2_inv_1_0.Y 0.00334f
C495 a_14538_17044# sg13g2_inv_1_0.Y 0.00345f
C496 sg13g2_a22oi_1_0.B2 a_15688_25154# 0
C497 sg13g2_dfrbpq_1_3.Q a_16735_16388# 0.01722f
C498 a_16266_15996# sg13g2_inv_1_1.A 0.0029f
C499 a_14248_23556# sg13g2_a21oi_1_0.A2 0.00763f
C500 sg13g2_inv_2_1.A sg13g2_inv_1_0.Y 0
C501 a_11940_14040# a_12817_14018# 0
C502 a_11654_13722# a_12297_14113# 0.00801f
C503 a_12357_13701# a_12459_13844# 0.47622f
C504 sg13g2_a22oi_1_0.B2 sg13g2_inv_1_0.Y 0.01117f
C505 a_14912_16668# VDD 0
C506 a_14061_12256# VDD 0.41908f
C507 a_16048_15454# a_15856_16238# 0
C508 a_15791_15311# a_15599_16357# 0.00198f
C509 a_15784_14570# sg13g2_dfrbpq_1_1.Q 0.00226f
C510 sg13g2_inv_1_0.Y a_12817_14018# 0.02121f
C511 a_12969_17137# sg13g2_a21oi_1_0.A2 0
C512 a_12459_13844# a_13456_13942# 0.02979f
C513 a_12652_16119# sg13g2_dfrbpq_1_0.CLK 0
C514 a_13864_16082# a_13131_16868# 0
C515 a_7816_15996# VDD 0.31209f
C516 a_25856_11890# VDD 0
C517 a_11493_16007# a_12134_14922# 0
C518 wake_up_sg a_11050_15964# 0
C519 sg13g2_dfrbpq_1_0.CLK a_12939_14495# 0.04495f
C520 a_14340_16000# sg13g2_dfrbpq_1_5.Q 0.00102f
C521 a_14697_16043# a_14314_15964# 0.00333f
C522 sg13g2_a21oi_1_0.A1 a_14054_16434# 0.01545f
C523 sg13g2_dfrbpq_1_3.D a_13679_14845# 0.0039f
C524 a_12612_17064# sg13g2_a21oi_1_0.A2 0.05704f
C525 a_13456_13942# a_13516_14037# 0.01042f
C526 a_15856_16238# sg13g2_dfrbpq_1_0.CLK 0.00322f
C527 a_13480_10620# VDD 0.0024f
C528 sg13g2_dfrbpq_1_0.CLK a_13297_14486# 0.00692f
C529 a_12592_16238# a_12394_14452# 0
C530 a_12900_16759# sg13g2_a21oi_1_0.A2 0
C531 a_11914_13945# a_11940_14040# 0.36952f
C532 sc_en VDD 0.33721f
C533 a_14532_14040# a_14346_14484# 0
C534 sg13g2_inv_1_0.Y a_11914_13945# 0.26965f
C535 a_15217_15998# VDD 0.0078f
C536 a_13664_10830# sg13g2_buf_1_4.A 0.0219f
C537 a_12652_16119# a_12335_16357# 0.00247f
C538 a_14248_23556# VDD 0.28393f
C539 Timer_en a_14144_4782# 0.00275f
C540 a_15791_13799# a_16294_14484# 0
C541 sg13g2_nor2_1_0.B a_12394_14452# 0.0039f
C542 a_14757_16007# sg13g2_dfrbpq_1_6.D 0.00214f
C543 a_14889_15625# VDD 0
C544 a_14061_12256# a_14155_12256# 0.00273f
C545 a_14757_16007# sg13g2_o21ai_1_0.A1 0.00431f
C546 a_13499_15996# sg13g2_nor2_1_0.B 0
C547 sg13g2_dfrbpq_1_4.D a_11050_15964# 0.01923f
C548 a_12969_17137# VDD 0
C549 a_15217_16349# sg13g2_dfrbpq_1_6.D 0.00171f
C550 sg13g2_dfrbpq_1_3.Q a_15791_13799# 0.00135f
C551 a_14506_15457# a_14054_16434# 0
C552 a_14532_15552# a_15784_14570# 0
C553 a_17800_15272# VDD 0.26811f
C554 sg13g2_inv_1_0.Y a_12420_14488# 0.43912f
C555 sg13g2_inv_1_1.A sg13g2_dfrbpq_1_1.Q 0.02284f
C556 a_13199_13799# a_12420_14488# 0
C557 sg13g2_a21oi_1_0.A1 sg13g2_inv_1_1.Y 0.01806f
C558 sg13g2_dfrbpq_1_4.D a_12592_16238# 0.00649f
C559 a_12459_13844# a_12939_14495# 0
C560 sg13g2_inv_1_1.A a_13996_14607# 0
C561 a_12612_17064# VDD 0.07873f
C562 sg13g2_a22oi_1_0.B2 a_14859_16007# 0.02629f
C563 a_15791_15311# a_15784_14570# 0
C564 a_16832_15366# VDD 0.0815f
C565 a_13864_16082# sg13g2_inv_1_0.Y 0
C566 a_15505_16357# a_15496_16878# 0
C567 a_12900_16759# VDD 0.00678f
C568 sg13g2_inv_1_0.Y a_13679_14845# 0.14653f
C569 a_12650_15532# VDD 0.00804f
C570 a_13401_14037# sg13g2_dfrbpq_1_0.CLK 0.00344f
C571 a_16048_15454# a_16051_14746# 0.00142f
C572 a_10024_15996# a_9920_16082# 0.00624f
C573 sg13g2_inv_1_1.A a_15801_16119# 0
C574 a_12357_13701# sg13g2_buf_1_0.A 0
C575 a_13199_13799# a_13679_14845# 0
C576 a_16458_15532# sg13g2_a21o_1_1.A2 0.00151f
C577 sg13g2_dfrbpq_1_4.D sg13g2_nor2_1_0.B 0.15506f
C578 a_16266_15996# sg13g2_inv_1_0.Y 0
C579 a_14235_17564# sg13g2_inv_1_0.Y 0
C580 a_14246_13722# VDD 0.80131f
C581 sg13g2_dfrbpq_1_5.Q VDD 0.57264f
C582 a_16210_15234# sg13g2_a21o_1_1.A2 0
C583 a_13456_13942# sg13g2_buf_1_0.A 0.00985f
C584 a_16210_13722# a_15791_13799# 0.00174f
C585 a_11364_16421# VDD 0.00601f
C586 sg13g2_dfrbpq_1_6.D a_14314_15964# 0
C587 sg13g2_dfrbpq_1_3.D sg13g2_dfrbpq_1_1.Q 0.00524f
C588 sg13g2_dfrbpq_1_0.CLK a_16051_14746# 0.00338f
C589 a_14757_16007# sg13g2_o21ai_1_0.B1 0
C590 a_14506_15457# sg13g2_inv_1_1.Y 0
C591 a_14340_13722# VDD 0
C592 a_12134_14922# a_12420_14488# 0.41329f
C593 a_12754_16434# VDD 0
C594 a_11848_15156# sg13g2_nor2_1_0.A 0.00241f
C595 adc_start a_16458_14020# 0
C596 sg13g2_a21oi_1_0.A1 a_15505_16357# 0
C597 timer_done a_13960_4782# 0
C598 a_14246_15234# a_14532_15552# 0.41329f
C599 a_16832_15366# a_16735_15972# 0
C600 a_14820_13735# VDD 0.0085f
C601 a_15217_16349# sg13g2_o21ai_1_0.B1 0
C602 a_14949_13701# sg13g2_dfrbpq_1_1.Q 0
C603 a_15051_13844# a_15784_14570# 0
C604 a_12228_13735# sg13g2_nor2_1_0.B 0
C605 a_14532_15552# sg13g2_inv_1_1.A 0.01632f
C606 a_15496_16878# sg13g2_dfrbpq_1_0.CLK 0.00121f
C607 a_13192_12342# sg13g2_dfrbpq_1_0.CLK 0
C608 a_14248_4688# a_14144_4782# 0.00624f
C609 sg13g2_nor2b_1_0.Y VDD 0.36901f
C610 a_12134_14922# a_13679_14845# 0
C611 a_12420_14488# a_13297_14837# 0.01835f
C612 a_12394_14452# a_12939_14495# 0.01f
C613 a_12837_14495# a_12708_14909# 0.01562f
C614 sg13g2_a21oi_1_0.A1 tx_start 0.19049f
C615 a_15872_25498# VDD 0
C616 a_15096_17064# a_14998_16742# 0.00202f
C617 a_14246_15234# a_15791_15311# 0
C618 a_16048_13942# sg13g2_dfrbpq_1_1.Q 0.00197f
C619 a_13401_14037# a_12459_13844# 0
C620 a_12166_13735# a_11940_14040# 0.0052f
C621 a_12228_13735# a_12357_13701# 0.01562f
C622 a_14340_16000# a_14628_16421# 0.43707f
C623 a_25856_17594# VDD 0.08554f
C624 a_15791_15311# sg13g2_inv_1_1.A 0.01731f
C625 a_13459_12404# VDD 0.33748f
C626 a_16735_15972# sg13g2_dfrbpq_1_5.Q 0.04761f
C627 a_12939_14495# a_13936_14726# 0.03061f
C628 a_11464_13644# VDD 0.00177f
C629 a_9920_16426# sg13g2_dfrbpq_1_0.CLK 0
C630 sg13g2_and2_1_0.X VDD 0.80231f
C631 a_12166_13735# sg13g2_inv_1_0.Y 0
C632 a_14532_15552# a_14820_15247# 0.43707f
C633 sg13g2_inv_1_1.A a_13871_16823# 0
C634 a_14340_16000# sg13g2_a21oi_1_0.A2 0.00165f
C635 a_13459_12404# a_13105_13799# 0
C636 sg13g2_buf_1_0.A a_13472_4782# 0.02359f
C637 sg13g2_buf_1_4.A a_14506_13945# 0
C638 a_14757_16007# sg13g2_dfrbpq_1_3.Q 0
C639 a_15697_13799# a_15784_14570# 0
C640 sg13g2_a21oi_1_0.A1 a_14128_16966# 0.0071f
C641 sg13g2_nor2_1_0.A a_10790_16434# 0.00393f
C642 a_14346_14484# a_14098_14922# 0
C643 a_14998_16742# sg13g2_dfrbpq_1_6.D 0.10668f
C644 sg13g2_buf_1_5.X a_14152_10736# 0.28141f
C645 a_17024_13644# sg13g2_a21o_1_1.A2 0
C646 a_16048_15454# a_15993_15549# 0.00412f
C647 sg13g2_o21ai_1_0.A1 a_14998_16742# 0.10047f
C648 a_14628_16421# sg13g2_a21oi_1_0.A2 0
C649 sg13g2_inv_1_0.Y sg13g2_dfrbpq_1_1.Q 0.00108f
C650 sg13g2_o21ai_1_0.B1 a_14314_15964# 0
C651 a_15856_16238# a_15599_16357# 0.34468f
C652 a_13585_14845# sg13g2_a21oi_1_0.A2 0
C653 sg13g2_dfrbpq_1_3.D a_14532_15552# 0.04268f
C654 a_14506_15457# a_14949_15213# 0.02242f
C655 a_12652_16119# sg13g2_dfrbpq_1_4.D 0
C656 sg13g2_inv_1_0.Y a_13996_14607# 0.01431f
C657 sg13g2_dfrbpq_1_4.D a_12939_14495# 0
C658 sg13g2_a21oi_1_0.A1 sg13g2_dfrbpq_1_0.CLK 0.57077f
C659 sg13g2_inv_1_1.A a_13777_16823# 0
C660 a_16018_16434# sg13g2_dfrbpq_1_5.Q 0
C661 sg13g2_a22oi_1_0.B2 a_14912_16668# 0.00112f
C662 sg13g2_a21oi_1_0.A1 a_14290_16746# 0
C663 a_11464_13854# VDD 0.15557f
C664 a_12592_16238# sg13g2_nor2_1_0.Y 0.04449f
C665 a_14152_10736# Timer_en 0.08749f
C666 a_16458_15532# a_16210_15234# 0
C667 a_14757_16007# a_14054_16434# 0.02432f
C668 a_14820_15247# a_14758_15247# 0
C669 a_14949_15213# a_14532_14040# 0
C670 a_15051_15356# sg13g2_dfrbpq_1_5.Q 0
C671 sg13g2_dfrbpq_1_3.D a_15791_15311# 0.01921f
C672 a_14532_15552# a_14949_13701# 0
C673 sg13g2_nor2_1_0.A a_11433_16043# 0
C674 a_15801_16119# sg13g2_inv_1_0.Y 0.00351f
C675 sg13g2_dfrbpq_1_0.CLK a_12136_16668# 0.00194f
C676 a_12817_13743# sg13g2_a21o_1_0.X 0.00118f
C677 sg13g2_a21oi_1_0.A1 a_11076_16000# 0
C678 a_13029_16725# a_14128_16966# 0
C679 a_13131_16868# a_13871_16823# 0.26905f
C680 sg13g2_dfrbpq_1_4.D a_13297_14486# 0
C681 a_17696_15366# VDD 0.09234f
C682 uart_en VDD 0.17827f
C683 a_25856_16878# a_25856_17594# 0
C684 a_15993_15549# sg13g2_dfrbpq_1_0.CLK 0
C685 a_14440_5412# Timer_en 0.00334f
C686 sg13g2_nor2_1_0.B sg13g2_nor2_1_0.Y 0.24938f
C687 a_13576_4688# VDD 0.26091f
C688 a_14155_12256# sg13g2_and2_1_0.X 0.00112f
C689 sg13g2_a21o_1_0.A2 a_13838_12256# 0
C690 a_14314_15964# a_14346_14484# 0
C691 sg13g2_dfrbpq_1_3.D a_14758_15247# 0
C692 sg13g2_nor2_1_0.A a_11654_13722# 0.00114f
C693 adc_en a_14144_4782# 0.00179f
C694 sg13g2_a21oi_1_0.A1 a_12335_16357# 0
C695 a_14340_16000# VDD 0.10215f
C696 a_13131_16868# a_13489_17042# 0.02138f
C697 a_13029_16725# sg13g2_dfrbpq_1_0.CLK 0.26754f
C698 sg13g2_inv_1_1.A a_16108_14037# 0
C699 sg13g2_inv_1_1.A adc_done 0.00169f
C700 a_14246_15234# sg13g2_nor2_1_0.B 0
C701 a_13459_12404# a_13480_10830# 0
C702 sg13g2_a21oi_1_0.A1 a_14188_17061# 0.00134f
C703 a_14506_15457# sg13g2_dfrbpq_1_0.CLK 0.00419f
C704 a_13960_4572# VDD 0.00206f
C705 a_12838_16759# sg13g2_dfrbpq_1_0.CLK 0
C706 a_13777_16823# a_13131_16868# 0.00647f
C707 a_25768_14570# VDD 0.15802f
C708 a_14148_16434# sg13g2_a21oi_1_0.A2 0
C709 a_15697_15311# sg13g2_dfrbpq_1_5.Q 0
C710 a_13866_14020# a_13679_14845# 0
C711 a_16048_15454# a_15791_13799# 0
C712 a_15791_15311# a_16048_13942# 0
C713 sg13g2_a21o_1_1.A2 a_16832_15156# 0.00232f
C714 sg13g2_inv_1_1.A sg13g2_nor2_1_0.B 0
C715 a_14628_16421# VDD 0.008f
C716 sg13g2_a22oi_1_0.B2 a_15217_15998# 0
C717 sg13g2_dfrbpq_1_0.CLK a_10790_16434# 0.0156f
C718 a_13585_14845# VDD 0.00479f
C719 sg13g2_a22oi_1_0.B2 a_14248_23556# 0
C720 tx_start a_15976_25068# 0
C721 a_12134_14922# a_13996_14607# 0
C722 a_14532_14040# sg13g2_dfrbpq_1_0.CLK 0.07449f
C723 a_14998_16742# sg13g2_o21ai_1_0.B1 0.03467f
C724 a_13401_14037# sg13g2_buf_1_0.A 0
C725 sg13g2_a21oi_1_0.A2 VDD 2.5718f
C726 a_14532_15552# sg13g2_inv_1_0.Y 0.4149f
C727 a_14757_16007# sg13g2_inv_1_1.Y 0
C728 a_16430_14832# a_16051_14746# 0
C729 sg13g2_dfrbpq_1_3.D a_15051_13844# 0.00277f
C730 a_16294_14484# sg13g2_a21o_1_1.A2 0.01685f
C731 sg13g2_dfrbpq_1_0.CLK a_11953_16349# 0.00332f
C732 a_13029_16725# a_12335_16357# 0.00312f
C733 a_12612_17064# a_13002_15996# 0
C734 a_10790_16434# a_11076_16000# 0.41329f
C735 sg13g2_dfrbpq_1_6.D a_12326_16746# 0.29362f
C736 a_17800_15272# sg13g2_inv_2_1.A 0.26119f
C737 a_15791_13799# sg13g2_dfrbpq_1_0.CLK 0.00372f
C738 a_12939_14495# a_13881_14607# 0
C739 a_14054_16434# a_14314_15964# 0.75507f
C740 a_15856_16238# a_15784_14570# 0
C741 a_15791_15311# sg13g2_inv_1_0.Y 0.13303f
C742 a_14073_17061# sg13g2_dfrbpq_1_6.D 0
C743 a_14532_14040# a_15409_14018# 0
C744 a_14246_13722# a_14889_14113# 0.00801f
C745 a_14949_13701# a_15051_13844# 0.47622f
C746 a_10790_16434# a_12335_16357# 0
C747 a_11050_15964# a_11595_16007# 0.01f
C748 a_11076_16000# a_11953_16349# 0.01835f
C749 a_11493_16007# a_11364_16421# 0.01562f
C750 sg13g2_nor2_1_0.A sg13g2_a21o_1_0.X 0
C751 sg13g2_inv_1_1.Y a_14098_14922# 0
C752 a_15599_16357# a_16051_14746# 0
C753 reset a_8776_13644# 0.00207f
C754 a_16832_15366# sg13g2_inv_2_1.A 0.019f
C755 sg13g2_inv_1_0.Y a_13871_16823# 0.14402f
C756 sg13g2_dfrbpq_1_3.D sg13g2_nor2_1_0.B 0
C757 sg13g2_dfrbpq_1_3.Q sg13g2_a21o_1_1.A2 0.30602f
C758 a_16832_15366# sg13g2_a22oi_1_0.B2 0
C759 a_15096_17064# sg13g2_dfrbpq_1_6.D 0.01075f
C760 a_14758_15247# sg13g2_inv_1_0.Y 0
C761 a_14148_16434# VDD 0
C762 a_13768_10736# timer_done 0.01199f
C763 sg13g2_dfrbpq_1_0.CLK a_11654_13722# 0
C764 a_15051_13844# a_16048_13942# 0.02979f
C765 a_14859_16007# a_15801_16119# 0
C766 a_11595_16007# a_12592_16238# 0.03061f
C767 sg13g2_dfrbpq_1_3.D a_15697_13799# 0
C768 sg13g2_o21ai_1_0.A1 a_15096_17064# 0.00139f
C769 a_12586_16969# sg13g2_dfrbpq_1_0.CLK 0
C770 sg13g2_inv_1_0.Y a_13489_17042# 0.01491f
C771 sg13g2_inv_2_1.A sg13g2_dfrbpq_1_5.Q 0.00612f
C772 a_13192_12342# sg13g2_buf_1_0.A 0.00152f
C773 sg13g2_nor2b_1_0.Y a_11493_16007# 0.00272f
C774 a_14336_5842# timer_done 0.00106f
C775 a_13777_16823# sg13g2_inv_1_0.Y 0
C776 sg13g2_a22oi_1_0.B2 sg13g2_dfrbpq_1_5.Q 0.3115f
C777 a_13002_15996# a_12754_16434# 0
C778 a_11595_16007# sg13g2_nor2_1_0.B 0
C779 a_16048_13942# a_16108_14037# 0.01042f
C780 a_15051_13844# a_15409_13743# 0.00104f
C781 a_14949_13701# a_15697_13799# 0.01058f
C782 a_15791_13799# a_16458_14020# 0.0894f
C783 a_14440_5412# a_14248_4688# 0
C784 a_12652_16119# sg13g2_nor2_1_0.Y 0
C785 a_14757_16007# a_15505_16357# 0.01058f
C786 sg13g2_nor2_1_0.Y a_12939_14495# 0
C787 sg13g2_dfrbpq_1_6.D a_12241_16357# 0.00206f
C788 sg13g2_inv_1_0.Y a_11050_15964# 0.2637f
C789 a_13105_13799# VDD 0.00294f
C790 a_16048_13942# a_15697_13799# 0.008f
C791 a_15051_13844# sg13g2_inv_1_0.Y 0.42489f
C792 sg13g2_inv_1_1.Y a_14314_15964# 0.00404f
C793 a_14949_15213# a_14757_16007# 0
C794 sg13g2_o21ai_1_0.A1 sg13g2_dfrbpq_1_6.D 0.34452f
C795 sg13g2_nor2b_1_0.Y a_12136_16878# 0
C796 sg13g2_nor2_1_0.Y a_13297_14486# 0
C797 a_11848_15366# sg13g2_nor2b_1_0.Y 0.00444f
C798 sg13g2_inv_1_0.Y a_12592_16238# 0.12835f
C799 a_12586_16969# a_12335_16357# 0
C800 sg13g2_a21oi_1_0.A1 a_13499_15996# 0.03306f
C801 sg13g2_a21oi_1_0.A1 a_13936_14726# 0
C802 uart_busy a_15872_25498# 0.00127f
C803 a_13664_10620# sg13g2_buf_1_0.A 0.00203f
C804 sg13g2_nor2_1_0.B a_11940_14040# 0
C805 a_14532_15552# a_14859_16007# 0
C806 a_16108_14037# sg13g2_inv_1_0.Y 0.01227f
C807 a_14144_23642# tx_start 0
C808 sg13g2_dfrbpq_1_0.CLK sg13g2_a21o_1_0.X 0.002f
C809 sg13g2_a22oi_1_0.B2 a_15872_25498# 0
C810 a_15856_16238# sg13g2_inv_1_1.A 0.00216f
C811 sg13g2_inv_1_0.Y sg13g2_nor2_1_0.B 0.26833f
C812 sg13g2_a21oi_1_0.A1 a_15599_16357# 0
C813 a_11654_13722# a_12459_13844# 0.097f
C814 a_11940_14040# a_12357_13701# 0.37291f
C815 sg13g2_buf_1_4.A sg13g2_inv_1_1.Y 0
C816 sg13g2_nor2_1_0.B a_13199_13799# 0
C817 a_15688_25154# a_15872_25154# 0.0524f
C818 a_15697_13799# sg13g2_inv_1_0.Y 0
C819 a_15096_17064# sg13g2_o21ai_1_0.B1 0
C820 a_13856_25498# VDD 0
C821 a_15784_14570# a_16051_14746# 0.00872f
C822 sg13g2_inv_1_0.Y a_12357_13701# 0.07392f
C823 a_16735_15972# VDD 0.30448f
C824 a_11654_13722# a_13516_14037# 0
C825 a_11940_14040# a_13456_13942# 0.00242f
C826 a_12357_13701# a_13199_13799# 0.00332f
C827 sg13g2_a21oi_1_0.A1 sg13g2_dfrbpq_1_4.D 0.11522f
C828 a_25856_16878# VDD 0.08554f
C829 a_14757_16007# sg13g2_dfrbpq_1_0.CLK 0.29738f
C830 a_13864_16082# a_12612_17064# 0
C831 a_14155_12256# VDD 0.00172f
C832 sg13g2_dfrbpq_1_0.CLK a_12708_14909# 0.0025f
C833 a_16458_15532# sg13g2_dfrbpq_1_3.Q 0.14438f
C834 a_14340_16000# a_14912_16878# 0
C835 wake_up_sg a_10790_16434# 0
C836 sg13g2_inv_1_0.Y a_13456_13942# 0.1139f
C837 a_14697_16043# a_14054_16434# 0.00801f
C838 clk a_7816_15996# 0.28839f
C839 a_13838_12256# sg13g2_buf_1_4.A 0.00232f
C840 a_13199_13799# a_13456_13942# 0.34468f
C841 a_15217_16349# sg13g2_dfrbpq_1_0.CLK 0.00105f
C842 sg13g2_nor2b_1_0.Y a_11914_13945# 0
C843 a_12592_16238# a_12134_14922# 0
C844 a_13480_10830# VDD 0.13808f
C845 sg13g2_dfrbpq_1_0.CLK a_14098_14922# 0
C846 sg13g2_o21ai_1_0.B1 sg13g2_dfrbpq_1_6.D 0.22379f
C847 a_16210_15234# sg13g2_dfrbpq_1_3.Q 0
C848 sg13g2_dfrbpq_1_3.D a_15856_16238# 0
C849 a_14246_13722# a_13679_14845# 0
C850 a_14152_10736# sg13g2_buf_1_4.A 0.00135f
C851 a_14506_15457# sg13g2_buf_1_0.A 0
C852 sg13g2_o21ai_1_0.A1 sg13g2_o21ai_1_0.B1 0.03551f
C853 a_16018_16434# VDD 0
C854 sg13g2_inv_1_0.Y a_8776_13644# 0
C855 a_25768_25154# VDD 0.13581f
C856 a_12537_16119# a_12592_16238# 0.00412f
C857 a_12652_16119# a_11595_16007# 0
C858 a_12335_16357# a_12708_14909# 0
C859 a_13029_16725# sg13g2_dfrbpq_1_4.D 0
C860 sg13g2_a21o_1_0.X a_12459_13844# 0.00127f
C861 a_14152_5498# VDD 0.1537f
C862 sg13g2_nor2_1_0.B a_12134_14922# 0.00347f
C863 Timer_en a_13472_4572# 0
C864 sg13g2_inv_2_1.A a_17696_15366# 0.00301f
C865 wake_up_sg a_11433_16043# 0
C866 a_16266_15996# sg13g2_dfrbpq_1_5.Q 0.12951f
C867 a_15051_15356# VDD 0.19201f
C868 a_14340_16000# a_14538_17044# 0
C869 a_14532_14040# sg13g2_buf_1_0.A 0.03105f
C870 sg13g2_buf_1_5.X sg13g2_buf_1_0.A 0.00377f
C871 a_15496_16878# a_15680_16878# 0.0524f
C872 sg13g2_nor2b_1_0.Y a_12420_14488# 0.00199f
C873 sg13g2_dfrbpq_1_4.D a_10790_16434# 0.28718f
C874 sg13g2_nor2_1_0.B a_13297_14837# 0
C875 a_14566_16421# sg13g2_dfrbpq_1_6.D 0
C876 sg13g2_a22oi_1_0.B2 a_14340_16000# 0.03762f
C877 a_16108_15549# VDD 0.00674f
C878 Timer_en sg13g2_buf_1_0.A 6.40005f
C879 a_14628_16421# a_14538_17044# 0
C880 sg13g2_inv_1_0.Y a_12228_14922# 0
C881 sg13g2_dfrbpq_1_0.CLK a_14314_15964# 0.0201f
C882 sg13g2_inv_1_1.A a_16051_14746# 0.00355f
C883 sg13g2_nor2_1_0.B a_12777_14531# 0
C884 sg13g2_a21oi_1_0.A1 a_13601_16344# 0.01147f
C885 a_12136_16878# sg13g2_a21oi_1_0.A2 0
C886 sg13g2_a22oi_1_0.B2 a_14628_16421# 0.00526f
C887 a_14538_17044# sg13g2_a21oi_1_0.A2 0.00231f
C888 a_15697_15311# VDD 0.0013f
C889 a_12652_16119# sg13g2_inv_1_0.Y 0.01938f
C890 sg13g2_inv_1_0.Y a_12939_14495# 0.43355f
C891 a_25672_11546# a_25856_11546# 0.0524f
C892 a_14506_13945# a_14346_14484# 0.00192f
C893 sg13g2_and2_1_0.X a_13679_14845# 0.00135f
C894 a_9920_16426# a_10024_15996# 0
C895 a_16048_15454# sg13g2_a21o_1_1.A2 0
C896 sg13g2_dfrbpq_1_4.D a_11433_16043# 0
C897 a_11654_13722# sg13g2_buf_1_0.A 0
C898 a_13199_13799# a_12939_14495# 0.00198f
C899 a_14949_15213# a_14998_16742# 0
C900 sg13g2_a22oi_1_0.B2 sg13g2_a21oi_1_0.A2 0.00121f
C901 a_15856_16238# sg13g2_inv_1_0.Y 0.09878f
C902 a_14912_16878# VDD 0.0765f
C903 sg13g2_inv_1_0.Y a_13297_14486# 0.01788f
C904 a_13768_10736# a_13480_10620# 0
C905 sg13g2_a21o_1_0.A2 sg13g2_buf_1_0.A 0.0051f
C906 sg13g2_buf_1_4.A sg13g2_dfrbpq_1_0.CLK 0.00113f
C907 a_11493_16007# VDD 0.2548f
C908 sg13g2_dfrbpq_1_6.D a_14054_16434# 0.00229f
C909 a_16832_15366# sg13g2_dfrbpq_1_1.Q 0
C910 a_14889_14113# VDD 0
C911 a_14073_17061# sg13g2_inv_1_1.Y 0
C912 sg13g2_dfrbpq_1_0.CLK sg13g2_a21o_1_1.A2 0
C913 sg13g2_dfrbpq_1_3.D a_16051_14746# 0.17615f
C914 a_12134_14922# a_12228_14922# 0.00716f
C915 adc_start a_16048_13942# 0
C916 a_13002_15996# VDD 0.38576f
C917 sg13g2_a21oi_1_0.A1 sg13g2_nor2_1_0.Y 0.03207f
C918 a_12136_16878# VDD 0.15258f
C919 a_14532_14040# a_15784_14570# 0
C920 a_14566_16421# sg13g2_o21ai_1_0.B1 0
C921 a_17128_13760# VDD 0.23761f
C922 a_14998_16742# sg13g2_dfrbpq_1_0.CLK 0.00111f
C923 a_14538_17044# VDD 0.38555f
C924 uart_busy VDD 0.1533f
C925 a_13576_4688# a_13960_4782# 0.01f
C926 a_14246_15234# sg13g2_a21oi_1_0.A1 0
C927 a_12394_14452# a_12708_14909# 0.00463f
C928 a_12420_14488# a_12646_14909# 0.0052f
C929 a_12134_14922# a_12939_14495# 0.097f
C930 a_11848_15366# VDD 0.16361f
C931 a_14144_23986# tx_start 0
C932 a_16735_16388# sg13g2_inv_1_1.A 0.00132f
C933 sg13g2_a21o_1_0.X sg13g2_buf_1_0.A 0.03538f
C934 sg13g2_inv_2_1.A VDD 0.83109f
C935 a_14437_17878# sg13g2_a21oi_1_0.A2 0
C936 a_14949_15213# a_15409_15530# 0.01483f
C937 sg13g2_a21oi_1_0.A1 sg13g2_inv_1_1.A 0
C938 sg13g2_nor2b_1_0.Y a_12166_13735# 0
C939 a_15791_13799# a_15784_14570# 0
C940 a_12228_13735# a_11654_13722# 0.31978f
C941 sg13g2_a22oi_1_0.B2 VDD 2.38189f
C942 sg13g2_dfrbpq_1_3.Q a_16832_15156# 0.00227f
C943 a_14340_16000# a_13679_14845# 0
C944 a_16840_13644# VDD 0.00177f
C945 a_15801_16119# sg13g2_dfrbpq_1_5.Q 0
C946 a_12817_14018# VDD 0.00761f
C947 a_12134_14922# a_13297_14486# 0
C948 a_12420_14488# a_13585_14845# 0.43239f
C949 a_13297_14837# a_12939_14495# 0.00104f
C950 a_16048_13942# a_16051_14746# 0.00138f
C951 a_16458_14020# sg13g2_a21o_1_1.A2 0.00125f
C952 sg13g2_buf_1_5.X a_13702_12532# 0
C953 a_13401_14037# sg13g2_inv_1_0.Y 0.00411f
C954 adc_start sg13g2_inv_1_0.Y 0
C955 sg13g2_dfrbpq_1_5.Q a_15496_16668# 0.0036f
C956 a_15051_15356# a_16108_15549# 0
C957 sg13g2_buf_1_0.A a_14248_4688# 0.27925f
C958 a_13029_16725# sg13g2_nor2_1_0.Y 0.0044f
C959 sg13g2_dfrbpq_1_6.D sg13g2_inv_1_1.Y 0
C960 a_12420_14488# sg13g2_a21oi_1_0.A2 0
C961 a_13866_14020# a_13456_13942# 0.10373f
C962 a_13401_14037# a_13199_13799# 0.00689f
C963 a_14757_16007# a_15599_16357# 0.00307f
C964 a_15993_15549# sg13g2_inv_1_1.A 0.00183f
C965 a_12838_16759# sg13g2_nor2_1_0.Y 0
C966 a_13864_16082# a_13585_14845# 0
C967 uart_done a_13856_25154# 0.02302f
C968 a_13679_14845# a_13585_14845# 0.28931f
C969 a_13936_14726# a_14098_14922# 0.00188f
C970 sg13g2_dfrbpq_1_3.Q a_16294_14484# 0.06804f
C971 a_10790_16434# sg13g2_nor2_1_0.Y 0
C972 a_15051_15356# a_15697_15311# 0.00647f
C973 sg13g2_buf_1_0.A a_14144_4572# 0
C974 a_13864_16082# sg13g2_a21oi_1_0.A2 0.01975f
C975 a_16048_15454# a_16458_15532# 0.10373f
C976 a_17024_13854# sg13g2_a21o_1_1.A2 0
C977 a_14859_16007# a_15856_16238# 0.03061f
C978 a_14697_16043# sg13g2_dfrbpq_1_0.CLK 0
C979 sg13g2_o21ai_1_0.B1 a_14054_16434# 0
C980 a_13679_14845# sg13g2_a21oi_1_0.A2 0
C981 a_14506_15457# a_14246_15234# 0.75507f
C982 a_14757_16007# sg13g2_dfrbpq_1_4.D 0
C983 sg13g2_a21oi_1_0.A1 a_13131_16868# 0.00109f
C984 a_14098_14922# sg13g2_buf_1_0.A 0
C985 sg13g2_inv_1_0.Y a_16051_14746# 0.00336f
C986 a_15916_16119# sg13g2_o21ai_1_0.A1 0
C987 a_14506_15457# sg13g2_inv_1_1.A 0.01954f
C988 a_15680_16668# sg13g2_dfrbpq_1_6.D 0
C989 sg13g2_a21oi_1_0.A1 a_13489_16767# 0
C990 a_11914_13945# VDD 0.09633f
C991 a_15409_15530# sg13g2_dfrbpq_1_0.CLK 0.00746f
C992 sg13g2_dfrbpq_1_3.D sg13g2_a21oi_1_0.A1 0
C993 a_13960_25068# sg13g2_a21oi_1_0.A2 0.27683f
C994 sg13g2_inv_2_1.A a_16735_15972# 0.03263f
C995 a_16048_15454# a_16210_15234# 0.00188f
C996 a_14235_17564# sg13g2_a21oi_1_0.A2 0.19758f
C997 a_14532_15552# sg13g2_dfrbpq_1_5.Q 0
C998 sg13g2_o21ai_1_0.A1 a_15680_16668# 0
C999 sg13g2_a22oi_1_0.B2 a_16735_15972# 0.06687f
C1000 a_12228_13735# sg13g2_a21o_1_0.X 0.00176f
C1001 sg13g2_nor2_1_0.A a_12241_16357# 0
C1002 a_14437_17878# VDD 0.00225f
C1003 a_12612_17064# a_13871_16823# 0.01529f
C1004 sg13g2_nor2_1_0.A sg13g2_dfrbpq_1_6.D 0
C1005 a_14073_17061# a_14128_16966# 0.00412f
C1006 a_16458_15532# sg13g2_dfrbpq_1_0.CLK 0.00102f
C1007 a_14152_5842# Timer_en 0.0043f
C1008 a_13192_12342# sg13g2_inv_1_0.Y 0
C1009 sg13g2_a21o_1_0.A2 a_13702_12532# 0.01543f
C1010 a_12268_15532# sg13g2_nor2_1_0.A 0
C1011 a_15791_15311# sg13g2_dfrbpq_1_5.Q 0.00206f
C1012 sg13g2_dfrbpq_1_3.D a_15993_15549# 0
C1013 a_14506_15457# a_14820_15247# 0.00463f
C1014 adc_en a_13472_4572# 0
C1015 sg13g2_a21oi_1_0.A1 a_11595_16007# 0
C1016 Timer_en a_14336_5498# 0.00186f
C1017 a_12420_14488# VDD 0.09197f
C1018 a_16840_13854# VDD 0.12896f
C1019 a_12612_17064# a_13489_17042# 0
C1020 a_12326_16746# sg13g2_dfrbpq_1_0.CLK 0.00266f
C1021 a_13029_16725# a_13131_16868# 0.47622f
C1022 sg13g2_inv_1_1.A a_15791_13799# 0
C1023 a_15505_16357# sg13g2_o21ai_1_0.A1 0.00156f
C1024 a_13960_4782# VDD 0.12486f
C1025 a_13777_16823# a_12612_17064# 0.43239f
C1026 a_13489_16767# a_13029_16725# 0.02396f
C1027 a_25768_14914# VDD 0.0025f
C1028 a_14949_15213# sg13g2_dfrbpq_1_6.D 0
C1029 a_13866_14020# a_12939_14495# 0
C1030 sg13g2_nor2_1_0.A a_12297_14113# 0
C1031 a_14949_15213# sg13g2_o21ai_1_0.A1 0
C1032 a_13864_16082# VDD 0.14373f
C1033 a_12586_16969# sg13g2_nor2_1_0.Y 0.00153f
C1034 a_13679_14845# VDD 0.20183f
C1035 a_14506_15457# sg13g2_dfrbpq_1_3.D 0.00465f
C1036 sg13g2_a22oi_1_0.B2 a_16018_16434# 0
C1037 tx_start a_15688_25498# 0
C1038 a_15051_15356# sg13g2_inv_2_1.A 0
C1039 adc_en sg13g2_buf_1_0.A 0.03686f
C1040 a_13960_25068# VDD 0.27901f
C1041 a_15051_15356# sg13g2_a22oi_1_0.B2 0.00172f
C1042 sg13g2_dfrbpq_1_4.D a_14314_15964# 0
C1043 a_17800_15272# adc_done 0.25767f
C1044 a_16458_15532# a_16458_14020# 0
C1045 a_14235_17564# VDD 0.29958f
C1046 a_10790_16434# a_10884_16434# 0.00716f
C1047 a_13702_12532# sg13g2_a21o_1_0.X 0
C1048 sg13g2_dfrbpq_1_3.D a_14532_14040# 0.00175f
C1049 a_16266_15996# VDD 0.38483f
C1050 sg13g2_dfrbpq_1_0.CLK a_11302_16421# 0
C1051 a_12612_17064# a_12592_16238# 0
C1052 a_12326_16746# a_12335_16357# 0
C1053 a_16430_14832# sg13g2_a21o_1_1.A2 0
C1054 sg13g2_a21oi_1_0.A1 sg13g2_inv_1_0.Y 0.01437f
C1055 sg13g2_dfrbpq_1_6.D a_14128_16966# 0.01201f
C1056 sg13g2_o21ai_1_0.A1 a_14128_16966# 0
C1057 a_14188_17061# a_12326_16746# 0
C1058 a_16108_15549# sg13g2_a22oi_1_0.B2 0.00104f
C1059 sg13g2_buf_1_4.A sg13g2_buf_1_0.A 2.89439f
C1060 a_11848_15156# sg13g2_inv_1_0.Y 0.0022f
C1061 a_14246_13722# a_15051_13844# 0.097f
C1062 a_14532_14040# a_14949_13701# 0.37291f
C1063 a_12612_17064# sg13g2_nor2_1_0.B 0
C1064 sg13g2_dfrbpq_1_0.CLK a_12241_16357# 0.00509f
C1065 a_11050_15964# a_11364_16421# 0.00463f
C1066 a_10790_16434# a_11595_16007# 0.097f
C1067 a_11076_16000# a_11302_16421# 0.0052f
C1068 sg13g2_dfrbpq_1_3.D a_15791_13799# 0
C1069 sg13g2_dfrbpq_1_6.D sg13g2_dfrbpq_1_0.CLK 0.14451f
C1070 sg13g2_inv_1_0.Y a_12136_16668# 0.00148f
C1071 a_12650_15532# sg13g2_nor2_1_0.B 0
C1072 a_15697_15311# sg13g2_inv_2_1.A 0
C1073 a_15993_14037# sg13g2_dfrbpq_1_0.CLK 0
C1074 a_14290_16746# sg13g2_dfrbpq_1_6.D 0
C1075 sg13g2_o21ai_1_0.A1 sg13g2_dfrbpq_1_0.CLK 0
C1076 a_13864_16426# sg13g2_a21oi_1_0.A2 0.00434f
C1077 a_15993_15549# sg13g2_inv_1_0.Y 0.00351f
C1078 a_14246_13722# a_16108_14037# 0
C1079 a_14532_14040# a_16048_13942# 0.00242f
C1080 a_14949_13701# a_15791_13799# 0.00332f
C1081 a_11953_16349# a_11595_16007# 0.00104f
C1082 a_11076_16000# a_12241_16357# 0.43239f
C1083 sg13g2_dfrbpq_1_3.D a_14758_13735# 0
C1084 a_10790_16434# a_11953_15998# 0
C1085 a_14538_17044# a_14912_16878# 0.01061f
C1086 a_12136_16878# a_11493_16007# 0
C1087 sg13g2_dfrbpq_1_6.D a_11076_16000# 0.0027f
C1088 sg13g2_inv_1_0.Y a_13029_16725# 0.03573f
C1089 a_12586_16969# a_13131_16868# 0.01f
C1090 a_13856_25498# a_13960_25068# 0
C1091 a_14506_13945# sg13g2_dfrbpq_1_0.CLK 0.00212f
C1092 sg13g2_a22oi_1_0.B2 a_14912_16878# 0.00118f
C1093 a_11848_15366# a_11493_16007# 0.0024f
C1094 a_12838_16759# sg13g2_inv_1_0.Y 0
C1095 a_14532_14040# a_15409_13743# 0.01835f
C1096 a_15051_13844# a_14820_13735# 0.12701f
C1097 a_15791_13799# a_16048_13942# 0.34468f
C1098 a_12592_16238# a_12754_16434# 0.00188f
C1099 a_12335_16357# a_12241_16357# 0.28931f
C1100 a_14506_15457# sg13g2_inv_1_0.Y 0.27187f
C1101 a_14949_15213# sg13g2_o21ai_1_0.B1 0
C1102 sg13g2_dfrbpq_1_3.Q a_15916_16119# 0
C1103 sg13g2_dfrbpq_1_6.D a_12335_16357# 0.00371f
C1104 sg13g2_nor2_1_0.Y a_12708_14909# 0
C1105 sg13g2_inv_1_0.Y a_10790_16434# 0.11209f
C1106 a_14336_5498# a_14248_4688# 0
C1107 a_12166_13735# VDD 0
C1108 clk VDD 0.65894f
C1109 sg13g2_buf_1_5.X sg13g2_inv_1_0.Y 0
C1110 sg13g2_inv_1_1.Y a_14054_16434# 0.26917f
C1111 a_14532_14040# sg13g2_inv_1_0.Y 0.38326f
C1112 a_14188_17061# sg13g2_dfrbpq_1_6.D 0.0018f
C1113 sg13g2_and2_1_0.X a_15051_13844# 0.00115f
C1114 uart_done tx_start 0.40981f
C1115 a_14757_16007# sg13g2_inv_1_1.A 0.00313f
C1116 reset a_8968_13760# 0.27187f
C1117 a_12046_15276# a_12268_15532# 0
C1118 sg13g2_inv_1_0.Y a_11953_16349# 0.00139f
C1119 sg13g2_inv_2_1.A a_17128_13760# 0
C1120 sg13g2_nor2b_1_0.Y sg13g2_nor2_1_0.B 0.19316f
C1121 a_13664_10830# sg13g2_buf_1_0.A 0.00635f
C1122 a_15791_13799# sg13g2_inv_1_0.Y 0.13309f
C1123 a_15916_16119# a_14054_16434# 0
C1124 a_13864_16426# VDD 0.0029f
C1125 sg13g2_a22oi_1_0.B2 uart_busy 0.01152f
C1126 sg13g2_dfrbpq_1_1.Q VDD 0.78964f
C1127 a_16840_13644# a_17128_13760# 0
C1128 a_16266_15996# a_16018_16434# 0
C1129 sg13g2_a22oi_1_0.B2 sg13g2_inv_2_1.A 0.20446f
C1130 sg13g2_inv_1_1.A a_14098_14922# 0
C1131 sg13g2_nor2b_1_0.Y a_12357_13701# 0
C1132 sg13g2_a21oi_1_0.A1 a_14859_16007# 0.00325f
C1133 a_14340_16000# a_13871_16823# 0.00213f
C1134 sg13g2_inv_1_0.Y a_11433_16043# 0
C1135 a_13996_14607# VDD 0.00816f
C1136 a_11654_13722# a_11940_14040# 0.41329f
C1137 tx_start a_13856_25154# 0
C1138 sg13g2_o21ai_1_0.B1 sg13g2_dfrbpq_1_0.CLK 0
C1139 a_14949_15213# sg13g2_dfrbpq_1_3.Q 0
C1140 a_15976_25068# a_15688_25154# 0.00536f
C1141 sg13g2_inv_1_0.Y a_11654_13722# 0.1326f
C1142 a_15801_16119# VDD 0
C1143 sg13g2_and2_1_0.X a_15697_13799# 0
C1144 a_14697_16043# sg13g2_dfrbpq_1_4.D 0
C1145 a_11654_13722# a_13199_13799# 0
C1146 a_13192_12132# VDD 0.00226f
C1147 a_16048_15454# sg13g2_dfrbpq_1_3.Q 0.00285f
C1148 a_15496_16668# VDD 0.00217f
C1149 a_12586_16969# sg13g2_inv_1_0.Y 0.2481f
C1150 sg13g2_dfrbpq_1_0.CLK a_12837_14495# 0.28366f
C1151 sg13g2_a21o_1_0.A2 sg13g2_inv_1_0.Y 0
C1152 sg13g2_dfrbpq_1_3.D a_14757_16007# 0
C1153 sg13g2_dfrbpq_1_0.CLK a_16294_14484# 0
C1154 sg13g2_buf_1_5.X timer_done 0.04183f
C1155 sg13g2_inv_1_0.Y a_11748_13722# 0
C1156 a_13871_16823# sg13g2_a21oi_1_0.A2 0.01596f
C1157 a_13702_12532# sg13g2_buf_1_4.A 0.08185f
C1158 a_13459_12404# a_13456_13942# 0
C1159 a_13768_10736# VDD 0.24991f
C1160 a_9920_16082# VDD 0.09231f
C1161 a_14246_15234# a_14314_15964# 0
C1162 sg13g2_dfrbpq_1_0.CLK a_14346_14484# 0.00188f
C1163 sg13g2_inv_1_1.A a_14314_15964# 0.00181f
C1164 a_16735_15972# sg13g2_dfrbpq_1_1.Q 0
C1165 a_13489_17042# sg13g2_a21oi_1_0.A2 0.00419f
C1166 timer_done Timer_en 2.27389f
C1167 adc_done a_17696_15366# 0.02303f
C1168 sg13g2_dfrbpq_1_3.Q sg13g2_dfrbpq_1_0.CLK 0.02791f
C1169 a_12335_16357# a_12837_14495# 0.00109f
C1170 sg13g2_a21o_1_0.X a_11940_14040# 0.00907f
C1171 a_14336_5842# VDD 0.00255f
C1172 a_13777_16823# sg13g2_a21oi_1_0.A2 0.0141f
C1173 a_15856_16238# sg13g2_dfrbpq_1_5.Q 0.0065f
C1174 a_14532_15552# VDD 0.09587f
C1175 a_16840_13854# a_17128_13760# 0.00536f
C1176 a_14128_16966# a_14054_16434# 0
C1177 sg13g2_nor2b_1_0.Y a_12228_14922# 0
C1178 sg13g2_inv_1_0.Y sg13g2_a21o_1_0.X 0.15319f
C1179 adc_done a_25768_14570# 0.00255f
C1180 sg13g2_a21o_1_0.X a_13199_13799# 0
C1181 a_15791_15311# VDD 0.17635f
C1182 sg13g2_inv_1_1.A sg13g2_buf_1_4.A 0
C1183 clk_gating_en sg13g2_buf_1_0.A 0.0021f
C1184 a_13618_13722# sg13g2_buf_1_0.A 0
C1185 sg13g2_dfrbpq_1_0.CLK a_14054_16434# 0.02387f
C1186 a_17800_15272# adc_start 0
C1187 a_12459_13844# a_12837_14495# 0
C1188 a_13871_16823# VDD 0.18863f
C1189 sg13g2_a22oi_1_0.B2 a_13864_16082# 0
C1190 a_14757_16007# sg13g2_inv_1_0.Y 0.0418f
C1191 sg13g2_inv_1_1.A sg13g2_a21o_1_1.A2 0.01042f
C1192 a_14758_15247# VDD 0
C1193 sg13g2_dfrbpq_1_3.Q a_16458_14020# 0
C1194 sg13g2_dfrbpq_1_3.D a_14314_15964# 0.00107f
C1195 a_14235_17564# a_14538_17044# 0
C1196 a_15599_16357# sg13g2_o21ai_1_0.A1 0.00137f
C1197 sg13g2_inv_1_0.Y a_12708_14909# 0.01117f
C1198 sg13g2_dfrbpq_1_4.D a_12241_16357# 0
C1199 sg13g2_inv_1_0.Y a_8968_13760# 0
C1200 a_13489_17042# VDD 0.00737f
C1201 sg13g2_a22oi_1_0.B2 a_14235_17564# 0
C1202 sg13g2_a22oi_1_0.B2 a_16266_15996# 0.01551f
C1203 sg13g2_dfrbpq_1_6.D sg13g2_dfrbpq_1_4.D 0
C1204 a_13777_16823# VDD 0.00374f
C1205 sg13g2_inv_1_0.Y a_14098_14922# 0
C1206 a_13768_10736# a_13480_10830# 0.00536f
C1207 sg13g2_a21oi_1_0.A1 a_14912_16668# 0.00305f
C1208 a_14144_17594# sg13g2_o21ai_1_0.B1 0
C1209 a_12817_13743# sg13g2_dfrbpq_1_0.CLK 0.00155f
C1210 a_12268_15532# sg13g2_dfrbpq_1_4.D 0
C1211 a_14506_13945# sg13g2_buf_1_0.A 0.03218f
C1212 a_14128_16966# sg13g2_inv_1_1.Y 0
C1213 a_11050_15964# VDD 0.10011f
C1214 a_8968_13760# a_8776_13854# 0.01209f
C1215 a_15051_13844# VDD 0.19677f
C1216 a_16210_13722# a_16458_14020# 0
C1217 a_12592_16238# VDD 0.16101f
C1218 sg13g2_dfrbpq_1_0.CLK sg13g2_inv_1_1.Y 0.08915f
C1219 sg13g2_dfrbpq_1_3.D sg13g2_a21o_1_1.A2 0.00223f
C1220 timer_done a_14248_4688# 0.04818f
C1221 a_16108_14037# VDD 0.00683f
C1222 adc_done VDD 1.70252f
C1223 a_14949_15213# a_15505_16357# 0
C1224 a_14248_4688# a_14632_4688# 0.0015f
C1225 a_13576_4688# a_13472_4782# 0.00624f
C1226 a_12134_14922# a_12708_14909# 0.31978f
C1227 a_12394_14452# a_12837_14495# 0.02242f
C1228 sg13g2_nor2_1_0.B VDD 0.61243f
C1229 a_14697_16043# sg13g2_inv_1_1.A 0
C1230 a_15916_16119# sg13g2_dfrbpq_1_0.CLK 0.00214f
C1231 a_14246_15234# a_15409_15530# 0
C1232 a_14532_15552# a_15051_15356# 0.34114f
C1233 sg13g2_inv_1_0.Y a_14314_15964# 0.26514f
C1234 timer_done a_14144_4572# 0.00139f
C1235 a_15697_13799# VDD 0.00289f
C1236 a_14248_23556# sg13g2_a21oi_1_0.A1 0.28481f
C1237 a_14235_17564# a_14437_17878# 0.01117f
C1238 a_13499_15996# a_12837_14495# 0
C1239 a_16430_14832# a_16294_14484# 0
C1240 a_15409_15530# sg13g2_inv_1_1.A 0.00263f
C1241 a_12420_14488# a_13679_14845# 0.01529f
C1242 a_12837_14495# a_13936_14726# 0
C1243 a_12708_14909# a_13297_14837# 0
C1244 a_12357_13701# VDD 0.25525f
C1245 a_15872_25154# VDD 0.06317f
C1246 sg13g2_buf_1_5.X a_14061_12256# 0.26753f
C1247 sg13g2_dfrbpq_1_5.Q a_15496_16878# 0.00376f
C1248 sg13g2_dfrbpq_1_6.D a_13601_16344# 0
C1249 a_12326_16746# sg13g2_nor2_1_0.Y 0.0022f
C1250 a_14949_15213# a_16048_15454# 0
C1251 a_15051_15356# a_15791_15311# 0.26905f
C1252 a_14340_16000# a_15856_16238# 0.00139f
C1253 a_14757_16007# a_14859_16007# 0.47795f
C1254 a_17128_13760# sg13g2_dfrbpq_1_1.Q 0.28934f
C1255 a_12817_13743# a_12459_13844# 0.00104f
C1256 a_13105_13799# a_12357_13701# 0.01058f
C1257 a_13864_16082# a_13679_14845# 0
C1258 a_16458_15532# sg13g2_inv_1_1.A 0.01694f
C1259 a_8968_13760# sg13g2_buf_1_6.X 0.24652f
C1260 sg13g2_nor2_1_0.A sg13g2_dfrbpq_1_0.CLK 0.04368f
C1261 a_12837_14495# sg13g2_buf_1_0.A 0
C1262 a_13936_14726# a_14346_14484# 0.10373f
C1263 a_12939_14495# a_13585_14845# 0.00647f
C1264 a_13456_13942# VDD 0.16565f
C1265 sg13g2_dfrbpq_1_3.Q a_16430_14832# 0.002f
C1266 sg13g2_inv_2_1.A sg13g2_dfrbpq_1_1.Q 0.01069f
C1267 sg13g2_buf_1_4.A sg13g2_inv_1_0.Y 0.02045f
C1268 a_15791_15311# a_16108_15549# 0.00247f
C1269 sg13g2_buf_1_0.A a_14144_4782# 0.02493f
C1270 a_14532_15552# a_15697_15311# 0.43239f
C1271 a_14949_15213# a_15409_15255# 0.02396f
C1272 sg13g2_a22oi_1_0.B2 sg13g2_dfrbpq_1_1.Q 0
C1273 sg13g2_buf_1_4.A a_13199_13799# 0.00147f
C1274 a_13105_13799# a_13456_13942# 0.008f
C1275 a_15217_16349# a_14859_16007# 0.00104f
C1276 a_12939_14495# sg13g2_a21oi_1_0.A2 0
C1277 a_15505_16357# sg13g2_dfrbpq_1_0.CLK 0.0023f
C1278 sg13g2_a21oi_1_0.A1 a_12612_17064# 0.00519f
C1279 a_16210_15234# sg13g2_inv_1_1.A 0
C1280 sg13g2_nor2_1_0.A a_11076_16000# 0.00133f
C1281 a_16840_13644# sg13g2_dfrbpq_1_1.Q 0.00624f
C1282 sg13g2_dfrbpq_1_4.D a_12837_14495# 0
C1283 a_14346_14484# sg13g2_buf_1_0.A 0.11665f
C1284 a_15680_16878# sg13g2_dfrbpq_1_6.D 0.00205f
C1285 sg13g2_inv_1_0.Y sg13g2_a21o_1_1.A2 0
C1286 a_14949_15213# sg13g2_dfrbpq_1_0.CLK 0.28261f
C1287 a_8776_13644# VDD 0.00177f
C1288 adc_done a_25856_16878# 0
C1289 a_15791_15311# a_15697_15311# 0.28931f
C1290 a_15599_16357# sg13g2_dfrbpq_1_3.Q 0.00253f
C1291 sg13g2_o21ai_1_0.A1 a_15680_16878# 0.00348f
C1292 sg13g2_a22oi_1_0.B2 a_15801_16119# 0
C1293 sg13g2_dfrbpq_1_3.D a_15409_15530# 0
C1294 a_14506_15457# a_14889_15625# 0.00333f
C1295 a_12326_16746# a_12420_16746# 0.00716f
C1296 sg13g2_nor2_1_0.A a_12335_16357# 0
C1297 a_16735_16388# sg13g2_dfrbpq_1_5.Q 0.00467f
C1298 a_16048_15454# sg13g2_dfrbpq_1_0.CLK 0.00164f
C1299 sg13g2_a22oi_1_0.B2 a_15496_16668# 0.00389f
C1300 a_14998_16742# sg13g2_inv_1_0.Y 0
C1301 sg13g2_a21oi_1_0.A1 sg13g2_dfrbpq_1_5.Q 0
C1302 sg13g2_a21o_1_0.A2 a_14061_12256# 0.00359f
C1303 a_13459_12404# a_13192_12342# 0.00872f
C1304 timer_done adc_en 0
C1305 a_15051_15356# a_15051_13844# 0
C1306 a_12046_15276# sg13g2_nor2_1_0.A 0.27095f
C1307 a_13499_15996# a_14054_16434# 0.00243f
C1308 sg13g2_dfrbpq_1_6.D sg13g2_nor2_1_0.Y 0.00217f
C1309 sg13g2_dfrbpq_1_3.D a_16458_15532# 0.00156f
C1310 sg13g2_dfrbpq_1_0.CLK a_14128_16966# 0
C1311 a_12228_14922# VDD 0
C1312 a_12612_17064# a_13029_16725# 0.37291f
C1313 a_12326_16746# a_13131_16868# 0.097f
C1314 a_15409_15255# sg13g2_dfrbpq_1_0.CLK 0.00635f
C1315 a_12268_15532# sg13g2_nor2_1_0.Y 0
C1316 a_14290_16746# a_14128_16966# 0.00188f
C1317 a_14073_17061# a_13131_16868# 0
C1318 a_12838_16759# a_12612_17064# 0.0052f
C1319 a_12900_16759# a_13029_16725# 0.01562f
C1320 a_13472_4782# VDD 0.07977f
C1321 a_15599_16357# a_14054_16434# 0
C1322 a_14859_16007# a_14314_15964# 0.01f
C1323 sg13g2_nor2_1_0.A a_12459_13844# 0
C1324 timer_done sg13g2_buf_1_4.A 0.00488f
C1325 sg13g2_a21oi_1_0.A1 a_12754_16434# 0
C1326 a_14246_15234# sg13g2_o21ai_1_0.A1 0
C1327 a_12652_16119# VDD 0.00648f
C1328 sg13g2_dfrbpq_1_3.D a_16210_15234# 0
C1329 a_12900_16759# a_12838_16759# 0
C1330 sg13g2_inv_1_1.A sg13g2_dfrbpq_1_6.D 0
C1331 adc_start a_25768_14570# 0.00173f
C1332 sg13g2_inv_1_1.A a_15993_14037# 0
C1333 a_12939_14495# VDD 0.20221f
C1334 sg13g2_inv_1_1.A sg13g2_o21ai_1_0.A1 0
C1335 a_14532_15552# sg13g2_inv_2_1.A 0
C1336 a_25768_4572# VDD 0.00121f
C1337 a_14532_15552# sg13g2_a22oi_1_0.B2 0
C1338 sg13g2_dfrbpq_1_4.D a_14054_16434# 0.00212f
C1339 a_15697_15311# a_15051_13844# 0
C1340 a_15856_16238# VDD 0.16243f
C1341 a_25768_23642# VDD 0.15447f
C1342 a_14061_12256# sg13g2_a21o_1_0.X 0
C1343 a_13297_14486# VDD 0.00826f
C1344 sg13g2_dfrbpq_1_0.CLK a_11076_16000# 0.10773f
C1345 a_12326_16746# a_11595_16007# 0
C1346 sg13g2_nor2b_1_0.Y a_11848_15156# 0.00418f
C1347 a_14697_16043# sg13g2_inv_1_0.Y 0
C1348 sg13g2_dfrbpq_1_6.D a_12420_16746# 0
C1349 a_16840_13854# sg13g2_dfrbpq_1_1.Q 0.03283f
C1350 a_15791_15311# sg13g2_inv_2_1.A 0.00212f
C1351 a_14188_17061# a_14128_16966# 0.01042f
C1352 a_14538_17044# a_13871_16823# 0.0894f
C1353 a_15409_14018# sg13g2_dfrbpq_1_0.CLK 0.00525f
C1354 a_15791_15311# sg13g2_a22oi_1_0.B2 0.00161f
C1355 a_12817_13743# sg13g2_buf_1_0.A 0
C1356 a_15409_15530# sg13g2_inv_1_0.Y 0.01621f
C1357 sg13g2_nor2b_1_0.Y a_12136_16668# 0
C1358 a_15680_16878# sg13g2_o21ai_1_0.B1 0
C1359 a_14820_15247# sg13g2_o21ai_1_0.A1 0
C1360 a_10790_16434# a_11364_16421# 0.31978f
C1361 a_11050_15964# a_11493_16007# 0.02242f
C1362 a_13499_15996# sg13g2_inv_1_1.Y 0.00659f
C1363 a_14246_13722# a_14532_14040# 0.41329f
C1364 sg13g2_dfrbpq_1_0.CLK a_12335_16357# 0.01736f
C1365 sg13g2_inv_1_1.Y a_13936_14726# 0
C1366 a_13679_14845# a_13996_14607# 0.00247f
C1367 a_12586_16969# a_12969_17137# 0.00333f
C1368 sg13g2_dfrbpq_1_6.D a_13131_16868# 0.02198f
C1369 a_14340_16000# a_15496_16878# 0
C1370 a_16458_14020# sg13g2_dfrbpq_1_0.CLK 0
C1371 sg13g2_o21ai_1_0.A1 a_13131_16868# 0
C1372 a_13489_16767# sg13g2_dfrbpq_1_6.D 0.00259f
C1373 a_16458_15532# sg13g2_inv_1_0.Y 0
C1374 a_16266_15996# sg13g2_dfrbpq_1_1.Q 0
C1375 sg13g2_dfrbpq_1_3.Q a_15784_14570# 0
C1376 a_12046_15276# sg13g2_dfrbpq_1_0.CLK 0
C1377 a_14246_13722# a_15791_13799# 0
C1378 a_11493_16007# a_12592_16238# 0
C1379 a_11364_16421# a_11953_16349# 0
C1380 a_11076_16000# a_12335_16357# 0.01529f
C1381 sg13g2_dfrbpq_1_3.D a_15993_14037# 0
C1382 sg13g2_inv_1_1.Y sg13g2_buf_1_0.A 0
C1383 sg13g2_dfrbpq_1_3.D sg13g2_o21ai_1_0.A1 0
C1384 sg13g2_inv_1_0.Y a_12326_16746# 0.08895f
C1385 a_12586_16969# a_12612_17064# 0.36952f
C1386 a_12046_15276# a_11076_16000# 0
C1387 sg13g2_nor2_1_0.A a_12394_14452# 0
C1388 a_17024_13854# sg13g2_dfrbpq_1_0.CLK 0
C1389 sg13g2_dfrbpq_1_0.CLK a_12459_13844# 0.03872f
C1390 a_12900_16759# a_12586_16969# 0.00463f
C1391 a_14073_17061# sg13g2_inv_1_0.Y 0.00351f
C1392 a_14532_14040# a_14820_13735# 0.43707f
C1393 wake_up_sg sg13g2_nor2_1_0.A 0.0276f
C1394 a_11493_16007# sg13g2_nor2_1_0.B 0.0019f
C1395 sg13g2_dfrbpq_1_4.D sg13g2_inv_1_1.Y 0
C1396 a_15599_16357# a_15916_16119# 0.00247f
C1397 a_12592_16238# a_13002_15996# 0.10373f
C1398 a_11595_16007# a_12241_16357# 0.00647f
C1399 sg13g2_dfrbpq_1_3.Q a_17006_16388# 0.00818f
C1400 sg13g2_dfrbpq_1_3.D a_14506_13945# 0.00131f
C1401 sc_en a_14248_4688# 0
C1402 sg13g2_nor2_1_0.Y a_12837_14495# 0
C1403 sg13g2_dfrbpq_1_6.D a_11595_16007# 0
C1404 sg13g2_inv_1_1.A sg13g2_o21ai_1_0.B1 0
C1405 sg13g2_inv_1_1.A a_16832_15156# 0
C1406 a_13401_14037# VDD 0
C1407 adc_start VDD 1.54847f
C1408 a_13838_12256# sg13g2_buf_1_0.A 0
C1409 sg13g2_dfrbpq_1_0.CLK a_13516_14037# 0.00414f
C1410 a_13002_15996# sg13g2_nor2_1_0.B 0.11615f
C1411 a_16048_13942# a_15993_14037# 0.00412f
C1412 sg13g2_buf_1_5.X sg13g2_and2_1_0.X 0.01806f
C1413 sg13g2_and2_1_0.X a_14532_14040# 0.05365f
C1414 a_14506_13945# a_14949_13701# 0.02242f
C1415 a_14757_16007# a_15217_15998# 0.01483f
C1416 sg13g2_inv_1_0.Y a_11302_16421# 0
C1417 a_12228_13735# a_12817_13743# 0
C1418 a_13866_14020# sg13g2_buf_1_4.A 0.12094f
C1419 sg13g2_a21oi_1_0.A1 a_14340_16000# 0.0382f
C1420 a_14144_17594# a_14128_16966# 0
C1421 sg13g2_inv_2_1.A adc_done 0.23942f
C1422 a_14152_10736# sg13g2_buf_1_0.A 0
C1423 a_14820_13735# a_14758_13735# 0
C1424 a_13618_13722# sg13g2_inv_1_0.Y 0
C1425 sg13g2_inv_1_1.A a_16294_14484# 0.00138f
C1426 sg13g2_and2_1_0.X a_15791_13799# 0
C1427 a_17800_15272# a_17696_15156# 0
C1428 a_13618_13722# a_13199_13799# 0.00174f
C1429 a_15856_16238# a_16018_16434# 0.00188f
C1430 a_15599_16357# a_15505_16357# 0.28931f
C1431 a_16051_14746# VDD 0.33625f
C1432 sg13g2_inv_1_0.Y a_12241_16357# 0.00979f
C1433 sg13g2_a21oi_1_0.A1 a_14628_16421# 0.01928f
C1434 a_14248_23556# a_14144_23642# 0.00624f
C1435 a_25768_25154# a_25768_23642# 0
C1436 sg13g2_nor2b_1_0.Y a_11654_13722# 0
C1437 uart_busy a_15872_25154# 0.02302f
C1438 sg13g2_nor2_1_0.B a_12817_14018# 0
C1439 sg13g2_nor2_1_0.A sg13g2_dfrbpq_1_4.D 0.11629f
C1440 a_14440_5412# sg13g2_buf_1_0.A 0.25844f
C1441 sg13g2_inv_1_0.Y sg13g2_dfrbpq_1_6.D 0.13773f
C1442 sg13g2_a21oi_1_0.A1 a_13585_14845# 0
C1443 a_15872_25498# a_15976_25068# 0
C1444 a_14949_15213# a_15599_16357# 0
C1445 a_15051_15356# a_15856_16238# 0
C1446 a_15993_14037# sg13g2_inv_1_0.Y 0.00351f
C1447 a_12268_15532# sg13g2_inv_1_0.Y 0
C1448 sg13g2_dfrbpq_1_3.D sg13g2_o21ai_1_0.B1 0
C1449 sg13g2_o21ai_1_0.A1 sg13g2_inv_1_0.Y 0
C1450 sg13g2_and2_1_0.X a_14758_13735# 0
C1451 sg13g2_dfrbpq_1_3.D a_16832_15156# 0
C1452 sg13g2_a22oi_1_0.B2 a_15872_25154# 0
C1453 sg13g2_dfrbpq_1_3.Q sg13g2_inv_1_1.A 0.48813f
C1454 sg13g2_a21oi_1_0.A1 sg13g2_a21oi_1_0.A2 0.93858f
C1455 a_13864_16082# a_13871_16823# 0
C1456 a_12357_13701# a_12817_14018# 0.01483f
C1457 a_11654_13722# a_11464_13644# 0.00404f
C1458 a_13192_12342# VDD 0.16299f
C1459 a_15496_16878# VDD 0.12716f
C1460 sg13g2_dfrbpq_1_0.CLK a_12394_14452# 0.00219f
C1461 a_16048_15454# a_15599_16357# 0.00123f
C1462 a_15791_15311# a_16266_15996# 0.00159f
C1463 wake_up_sg sg13g2_dfrbpq_1_0.CLK 0.34463f
C1464 a_13601_16344# sg13g2_inv_1_1.Y 0
C1465 a_14506_13945# sg13g2_inv_1_0.Y 0.26528f
C1466 a_13459_12404# sg13g2_a21o_1_0.A2 0.00148f
C1467 sg13g2_inv_1_0.Y a_12297_14113# 0.00108f
C1468 a_14061_12256# sg13g2_buf_1_4.A 0.16354f
C1469 a_12459_13844# a_13516_14037# 0
C1470 a_13499_15996# sg13g2_dfrbpq_1_0.CLK 0.0344f
C1471 a_14235_17564# a_13871_16823# 0.00163f
C1472 sg13g2_dfrbpq_1_0.CLK a_13936_14726# 0.00361f
C1473 a_9920_16426# VDD 0
C1474 a_25672_11546# VDD 0.13452f
C1475 a_13864_16082# a_13777_16823# 0
C1476 wake_up_sg a_11076_16000# 0
C1477 a_14757_16007# sg13g2_dfrbpq_1_5.Q 0
C1478 a_15697_15311# a_15856_16238# 0
C1479 sg13g2_nor2_1_0.B a_11914_13945# 0
C1480 sg13g2_dfrbpq_1_3.D a_14346_14484# 0.00532f
C1481 sg13g2_inv_1_1.A a_14054_16434# 0.00301f
C1482 Timer_en uart_en 0.00128f
C1483 a_12228_13735# sg13g2_nor2_1_0.A 0
C1484 sg13g2_a21oi_1_0.A1 a_14148_16434# 0
C1485 a_13029_16725# sg13g2_a21oi_1_0.A2 0.03181f
C1486 Timer_en a_13576_4688# 0.00441f
C1487 clk_gating_en a_14632_4688# 0.24489f
C1488 a_15599_16357# sg13g2_dfrbpq_1_0.CLK 0.0066f
C1489 a_13664_10620# VDD 0
C1490 a_12592_16238# a_12420_14488# 0
C1491 a_12335_16357# a_12394_14452# 0
C1492 a_11464_13854# a_11654_13722# 0.00201f
C1493 a_11914_13945# a_12357_13701# 0.02242f
C1494 sg13g2_dfrbpq_1_0.CLK sg13g2_buf_1_0.A 0.0292f
C1495 a_15217_16349# sg13g2_dfrbpq_1_5.Q 0
C1496 sg13g2_dfrbpq_1_3.D sg13g2_dfrbpq_1_3.Q 0.05039f
C1497 a_16735_16388# VDD 0
C1498 a_14998_16742# a_14912_16668# 0.00206f
C1499 sg13g2_inv_1_0.Y a_9728_13644# 0
C1500 a_13459_12404# sg13g2_a21o_1_0.X 0.18127f
C1501 sg13g2_nor2_1_0.B a_12420_14488# 0.00895f
C1502 Timer_en a_13960_4572# 0.00685f
C1503 sg13g2_a21oi_1_0.A1 VDD 2.24173f
C1504 sg13g2_dfrbpq_1_0.CLK sg13g2_dfrbpq_1_4.D 0.91997f
C1505 sg13g2_a21o_1_0.X a_11464_13644# 0.00444f
C1506 sg13g2_and2_1_0.X sg13g2_a21o_1_0.X 0
C1507 adc_done a_25768_14914# 0.00188f
C1508 a_11848_15156# VDD 0.00181f
C1509 sg13g2_o21ai_1_0.B1 sg13g2_inv_1_0.Y 0.00118f
C1510 a_15505_16357# a_15784_14570# 0
C1511 a_13702_12532# a_13838_12256# 0
C1512 sg13g2_dfrbpq_1_4.D a_11076_16000# 0.0185f
C1513 a_11940_14040# a_12837_14495# 0
C1514 a_13131_16868# a_14054_16434# 0
C1515 a_12136_16668# VDD 0.00121f
C1516 a_14859_16007# sg13g2_dfrbpq_1_6.D 0.00263f
C1517 a_14949_15213# a_15784_14570# 0.00104f
C1518 a_14246_15234# sg13g2_inv_1_1.Y 0.02997f
C1519 sg13g2_dfrbpq_1_3.D a_14054_16434# 0
C1520 a_15993_15549# VDD 0
C1521 a_14859_16007# sg13g2_o21ai_1_0.A1 0
C1522 sg13g2_inv_1_0.Y a_12837_14495# 0.04713f
C1523 sg13g2_inv_1_1.A sg13g2_inv_1_1.Y 0.11473f
C1524 a_13456_13942# a_12420_14488# 0
C1525 a_13199_13799# a_12837_14495# 0.00173f
C1526 sg13g2_dfrbpq_1_4.D a_12335_16357# 0.00886f
C1527 a_13029_16725# VDD 0.23908f
C1528 sg13g2_a22oi_1_0.B2 a_15856_16238# 0.01305f
C1529 a_15791_15311# sg13g2_dfrbpq_1_1.Q 0.00254f
C1530 a_14566_16421# sg13g2_inv_1_0.Y 0
C1531 a_11464_13854# sg13g2_a21o_1_0.X 0.03327f
C1532 a_14340_15234# sg13g2_inv_1_1.Y 0
C1533 a_15505_16357# a_15680_16878# 0
C1534 sg13g2_inv_1_0.Y a_14346_14484# 0.01923f
C1535 a_14506_15457# VDD 0.09995f
C1536 a_12838_16759# VDD 0
C1537 a_12228_13735# sg13g2_dfrbpq_1_0.CLK 0
C1538 a_12046_15276# sg13g2_dfrbpq_1_4.D 0.00173f
C1539 a_10024_15996# sg13g2_nor2_1_0.A 0.24593f
C1540 a_17800_15272# sg13g2_a21o_1_1.A2 0.00112f
C1541 a_12459_13844# sg13g2_buf_1_0.A 0
C1542 sg13g2_inv_1_1.A a_15916_16119# 0.00137f
C1543 a_16735_16388# a_16735_15972# 0
C1544 a_10790_16434# VDD 0.78695f
C1545 a_12586_16969# sg13g2_a21oi_1_0.A2 0.00171f
C1546 sg13g2_dfrbpq_1_3.Q sg13g2_inv_1_0.Y 0.00177f
C1547 sg13g2_nor2_1_0.A sg13g2_nor2_1_0.Y 0.0898f
C1548 sg13g2_buf_1_5.X VDD 0.94285f
C1549 a_14532_14040# VDD 0.09642f
C1550 a_15697_15311# a_16051_14746# 0
C1551 a_16832_15366# sg13g2_a21o_1_1.A2 0.00285f
C1552 a_13516_14037# sg13g2_buf_1_0.A 0
C1553 sg13g2_dfrbpq_1_0.CLK a_15784_14570# 0.00697f
C1554 a_11953_16349# VDD 0
C1555 a_16210_13722# a_16048_13942# 0.00188f
C1556 a_13866_14020# a_13618_13722# 0
C1557 sg13g2_buf_1_4.A a_14246_13722# 0.03688f
C1558 sg13g2_dfrbpq_1_0.CLK a_13601_16344# 0.00152f
C1559 a_13131_16868# sg13g2_inv_1_1.Y 0
C1560 sg13g2_inv_1_1.A sg13g2_nor2_1_0.A 0.00111f
C1561 uart_en a_14248_4688# 0.24499f
C1562 sg13g2_dfrbpq_1_0.CLK a_13881_14607# 0.00108f
C1563 a_15791_13799# VDD 0.18497f
C1564 sg13g2_buf_1_6.X a_9728_13644# 0.00121f
C1565 a_14152_5842# a_14440_5412# 0
C1566 Timer_en VDD 0.94498f
C1567 sg13g2_dfrbpq_1_3.D sg13g2_inv_1_1.Y 0.05216f
C1568 a_13576_4688# a_14248_4688# 0
C1569 a_12134_14922# a_12837_14495# 0.02432f
C1570 adc_start a_17128_13760# 0.24584f
C1571 a_11433_16043# VDD 0
C1572 sg13g2_dfrbpq_1_5.Q sg13g2_a21o_1_1.A2 0.00349f
C1573 sg13g2_buf_1_4.A a_14340_13722# 0
C1574 sg13g2_inv_1_0.Y a_14054_16434# 0.12637f
C1575 a_14440_5412# a_14336_5498# 0.00617f
C1576 a_14246_15234# a_14949_15213# 0.02454f
C1577 timer_done a_14144_4782# 0.00116f
C1578 sg13g2_a21oi_1_0.A1 a_16018_16434# 0
C1579 a_14758_13735# VDD 0
C1580 a_14144_23986# a_14248_23556# 0
C1581 a_14859_16007# sg13g2_o21ai_1_0.B1 0
C1582 a_14340_16000# a_14757_16007# 0.37384f
C1583 a_15051_13844# sg13g2_dfrbpq_1_1.Q 0
C1584 a_14248_4688# a_13960_4572# 0
C1585 a_14949_15213# sg13g2_inv_1_1.A 0.01628f
C1586 sg13g2_inv_2_1.A adc_start 0
C1587 a_12646_14909# a_12708_14909# 0
C1588 a_12837_14495# a_13297_14837# 0.02396f
C1589 a_12420_14488# a_12939_14495# 0.34102f
C1590 a_11654_13722# VDD 0.78247f
C1591 a_15976_25068# VDD 0.24955f
C1592 sg13g2_dfrbpq_1_5.Q a_14998_16742# 0
C1593 a_14532_15552# a_15791_15311# 0.01529f
C1594 a_16840_13644# adc_start 0.00192f
C1595 a_16108_14037# sg13g2_dfrbpq_1_1.Q 0
C1596 a_12817_13743# a_11940_14040# 0.01835f
C1597 a_12228_13735# a_12459_13844# 0.12701f
C1598 a_13866_14020# a_14506_13945# 0
C1599 a_14340_16000# a_15217_16349# 0.01835f
C1600 a_14757_16007# a_14628_16421# 0.01562f
C1601 a_12586_16969# VDD 0.09717f
C1602 sg13g2_a21o_1_0.A2 VDD 0.44683f
C1603 a_16048_15454# sg13g2_inv_1_1.A 0.0143f
C1604 a_13864_16082# a_12939_14495# 0
C1605 a_11748_13722# VDD 0
C1606 a_10024_15996# sg13g2_dfrbpq_1_0.CLK 0.01283f
C1607 a_12420_14488# a_13297_14486# 0
C1608 a_12939_14495# a_13679_14845# 0.26905f
C1609 sg13g2_buf_1_5.X a_14155_12256# 0.01071f
C1610 a_12817_13743# sg13g2_inv_1_0.Y 0.00227f
C1611 a_14532_15552# a_14758_15247# 0.0052f
C1612 sg13g2_inv_1_1.A a_14128_16966# 0
C1613 a_15051_15356# a_15993_15549# 0
C1614 a_14949_15213# a_14820_15247# 0.01562f
C1615 a_14757_16007# sg13g2_a21oi_1_0.A2 0
C1616 a_13459_12404# sg13g2_buf_1_4.A 0.01282f
C1617 sg13g2_buf_1_4.A sg13g2_and2_1_0.X 0.15615f
C1618 sg13g2_dfrbpq_1_0.CLK sg13g2_nor2_1_0.Y 0.14088f
C1619 a_14628_16421# a_15217_16349# 0
C1620 sg13g2_a22oi_1_0.B2 a_16051_14746# 0
C1621 a_15409_15255# sg13g2_inv_1_1.A 0
C1622 a_13585_14845# a_14098_14922# 0
C1623 a_13936_14726# sg13g2_buf_1_0.A 0.00128f
C1624 wake_up_sg sg13g2_dfrbpq_1_4.D 0.00922f
C1625 a_14246_15234# sg13g2_dfrbpq_1_0.CLK 0.00826f
C1626 a_14912_16668# sg13g2_dfrbpq_1_6.D 0
C1627 a_14144_23642# sg13g2_a21oi_1_0.A2 0.00338f
C1628 a_16458_15532# a_17800_15272# 0
C1629 sg13g2_inv_1_0.Y sg13g2_inv_1_1.Y 0.11018f
C1630 a_14859_16007# sg13g2_dfrbpq_1_3.Q 0
C1631 a_15856_16238# a_16266_15996# 0.10373f
C1632 sg13g2_inv_1_1.A sg13g2_dfrbpq_1_0.CLK 0.115f
C1633 sg13g2_dfrbpq_1_3.D a_14949_15213# 0.01365f
C1634 a_14506_15457# a_15051_15356# 0.01f
C1635 a_13499_15996# sg13g2_dfrbpq_1_4.D 0.15756f
C1636 sg13g2_nor2_1_0.A a_11595_16007# 0.00277f
C1637 a_12326_16746# a_12969_17137# 0.00801f
C1638 sg13g2_a21o_1_0.X VDD 0.97223f
C1639 sg13g2_a21oi_1_0.A1 a_14912_16878# 0.01629f
C1640 a_14340_15234# sg13g2_dfrbpq_1_0.CLK 0
C1641 sg13g2_a22oi_1_0.B2 a_15496_16878# 0.00165f
C1642 a_12335_16357# sg13g2_nor2_1_0.Y 0.02444f
C1643 a_14820_15247# a_15409_15255# 0
C1644 a_14340_16000# a_14314_15964# 0.36952f
C1645 sc_en clk_gating_en 4.07324f
C1646 a_16458_15532# a_16832_15366# 0.01061f
C1647 sg13g2_dfrbpq_1_3.D a_16048_15454# 0.00678f
C1648 a_14532_15552# a_15051_13844# 0
C1649 a_14949_15213# a_14949_13701# 0.00237f
C1650 sg13g2_nor2_1_0.A a_11953_15998# 0.00112f
C1651 a_15916_16119# sg13g2_inv_1_0.Y 0.01227f
C1652 sg13g2_dfrbpq_1_0.CLK a_12420_16746# 0
C1653 adc_en a_13576_4688# 0.24499f
C1654 a_13105_13799# sg13g2_a21o_1_0.X 0
C1655 sg13g2_a21oi_1_0.A1 a_11493_16007# 0
C1656 a_13131_16868# a_14128_16966# 0.02979f
C1657 a_12326_16746# a_12612_17064# 0.41329f
C1658 a_17696_15156# VDD 0
C1659 a_14820_15247# sg13g2_dfrbpq_1_0.CLK 0.00273f
C1660 a_13777_16823# a_13871_16823# 0.28931f
C1661 a_13838_12256# sg13g2_inv_1_0.Y 0
C1662 a_12900_16759# a_12326_16746# 0.31978f
C1663 a_14248_4688# VDD 0.25323f
C1664 sg13g2_a21o_1_0.A2 a_14155_12256# 0
C1665 a_14152_5498# Timer_en 0.00952f
C1666 a_16458_15532# sg13g2_dfrbpq_1_5.Q 0
C1667 a_14628_16421# a_14314_15964# 0.00463f
C1668 a_14859_16007# a_14054_16434# 0.097f
C1669 a_15791_15311# a_15051_13844# 0
C1670 a_15051_15356# a_15791_13799# 0
C1671 sg13g2_dfrbpq_1_3.D a_15409_15255# 0.0028f
C1672 sg13g2_nor2_1_0.A a_11940_14040# 0
C1673 sg13g2_a21oi_1_0.A1 a_13002_15996# 0
C1674 a_14757_16007# VDD 0.23714f
C1675 adc_en a_13960_4572# 0.00616f
C1676 adc_start a_25768_14914# 0
C1677 a_12708_14909# VDD 0.00957f
C1678 a_13131_16868# sg13g2_dfrbpq_1_0.CLK 0.0152f
C1679 a_14532_15552# sg13g2_nor2_1_0.B 0
C1680 a_14314_15964# sg13g2_a21oi_1_0.A2 0
C1681 sg13g2_nor2_1_0.A sg13g2_inv_1_0.Y 0.23317f
C1682 sg13g2_dfrbpq_1_3.D sg13g2_dfrbpq_1_0.CLK 0.08756f
C1683 a_8968_13760# VDD 0.25079f
C1684 a_14144_4572# VDD 0.00218f
C1685 a_13489_16767# sg13g2_dfrbpq_1_0.CLK 0.00932f
C1686 sg13g2_a21oi_1_0.A1 a_14538_17044# 0.14109f
C1687 a_16048_15454# a_16048_13942# 0
C1688 sg13g2_a21o_1_1.A2 a_17696_15366# 0
C1689 a_15217_16349# VDD 0.0014f
C1690 sg13g2_a22oi_1_0.B2 a_16735_16388# 0
C1691 sg13g2_dfrbpq_1_0.CLK a_10884_16434# 0
C1692 a_14144_23642# VDD 0.08585f
C1693 tx_start a_15688_25154# 0.00116f
C1694 a_15505_16357# sg13g2_inv_1_0.Y 0
C1695 sg13g2_dfrbpq_1_6.D a_12969_17137# 0
C1696 a_14098_14922# VDD 0
C1697 sg13g2_a22oi_1_0.B2 sg13g2_a21oi_1_0.A1 0.59937f
C1698 a_14949_13701# sg13g2_dfrbpq_1_0.CLK 0.27492f
C1699 a_12228_13735# sg13g2_buf_1_0.A 0
C1700 a_14949_15213# sg13g2_inv_1_0.Y 0.03847f
C1701 a_13499_15996# a_13601_16344# 0
C1702 a_13029_16725# a_13002_15996# 0.00351f
C1703 sg13g2_dfrbpq_1_0.CLK a_11595_16007# 0.03079f
C1704 a_10790_16434# a_11493_16007# 0.02432f
C1705 sg13g2_dfrbpq_1_3.D a_15409_14018# 0
C1706 sg13g2_dfrbpq_1_6.D a_12612_17064# 0.03855f
C1707 a_16048_13942# sg13g2_dfrbpq_1_0.CLK 0.00169f
C1708 a_13936_14726# a_13881_14607# 0.00412f
C1709 a_12939_14495# a_13996_14607# 0
C1710 a_12900_16759# sg13g2_dfrbpq_1_6.D 0.00768f
C1711 a_14188_17061# a_13131_16868# 0
C1712 sg13g2_o21ai_1_0.A1 a_12612_17064# 0
C1713 a_15993_15549# sg13g2_a22oi_1_0.B2 0
C1714 sg13g2_nor2b_1_0.Y a_12326_16746# 0
C1715 a_16048_15454# sg13g2_inv_1_0.Y 0.10177f
C1716 a_15599_16357# a_15784_14570# 0
C1717 a_11302_16421# a_11364_16421# 0
C1718 a_11493_16007# a_11953_16349# 0.02396f
C1719 a_11076_16000# a_11595_16007# 0.34102f
C1720 a_14859_16007# sg13g2_inv_1_1.Y 0
C1721 a_14949_13701# a_15409_14018# 0.01483f
C1722 a_13480_10830# sg13g2_a21o_1_0.X 0
C1723 sg13g2_dfrbpq_1_0.CLK a_11953_15998# 0
C1724 reset a_9728_13854# 0
C1725 sg13g2_inv_1_0.Y a_14128_16966# 0.10284f
C1726 sg13g2_buf_1_0.A a_13881_14607# 0
C1727 a_15409_13743# sg13g2_dfrbpq_1_0.CLK 0.00116f
C1728 sg13g2_dfrbpq_1_5.Q sg13g2_dfrbpq_1_6.D 0.02139f
C1729 a_15409_15255# sg13g2_inv_1_0.Y 0.00111f
C1730 sg13g2_nor2_1_0.A a_12134_14922# 0.002f
C1731 a_14152_10736# timer_done 0.26916f
C1732 a_14314_15964# VDD 0.11474f
C1733 sg13g2_dfrbpq_1_0.CLK a_11940_14040# 0.10394f
C1734 a_15051_13844# a_16108_14037# 0
C1735 sg13g2_dfrbpq_1_4.D a_13601_16344# 0.00663f
C1736 a_15856_16238# a_15801_16119# 0.00412f
C1737 a_14859_16007# a_15916_16119# 0
C1738 a_11595_16007# a_12335_16357# 0.26905f
C1739 wake_up_sg a_10024_15996# 0.26381f
C1740 a_11076_16000# a_11953_15998# 0
C1741 sg13g2_o21ai_1_0.A1 sg13g2_dfrbpq_1_5.Q 0.18261f
C1742 sg13g2_nor2_1_0.Y a_12394_14452# 0
C1743 a_15217_15998# sg13g2_o21ai_1_0.B1 0
C1744 sg13g2_inv_1_0.Y sg13g2_dfrbpq_1_0.CLK 0.58539f
C1745 a_15599_16357# a_15680_16878# 0
C1746 sg13g2_a21oi_1_0.A1 a_14437_17878# 0.00526f
C1747 a_12537_16119# sg13g2_nor2_1_0.A 0
C1748 adc_en VDD 0.14946f
C1749 a_12046_15276# a_11595_16007# 0
C1750 a_13702_12532# sg13g2_buf_1_0.A 0.09708f
C1751 sg13g2_dfrbpq_1_0.CLK a_13199_13799# 0.05264f
C1752 a_16048_13942# a_16458_14020# 0.10373f
C1753 a_15051_13844# a_15697_13799# 0.00647f
C1754 a_14440_5412# timer_done 0.05144f
C1755 a_12592_16238# sg13g2_nor2_1_0.B 0
C1756 a_12241_16357# a_12754_16434# 0
C1757 a_13499_15996# sg13g2_nor2_1_0.Y 0.00414f
C1758 a_14506_13945# a_14246_13722# 0.75507f
C1759 a_14440_5412# a_14632_4688# 0
C1760 a_14152_5498# a_14248_4688# 0
C1761 sg13g2_dfrbpq_1_6.D a_12754_16434# 0
C1762 sg13g2_inv_1_0.Y a_11076_16000# 0.38728f
C1763 sg13g2_a21oi_1_0.A1 a_12420_14488# 0
C1764 sg13g2_buf_1_4.A VDD 0.91842f
C1765 sg13g2_nor2b_1_0.Y a_12241_16357# 0
C1766 sg13g2_inv_1_1.A a_16430_14832# 0
C1767 a_15051_15356# a_14757_16007# 0
C1768 a_15409_14018# sg13g2_inv_1_0.Y 0.01621f
C1769 sg13g2_nor2b_1_0.Y sg13g2_dfrbpq_1_6.D 0.00172f
C1770 a_14859_16007# a_15505_16357# 0.00647f
C1771 sg13g2_inv_1_0.Y a_12335_16357# 0.16804f
C1772 a_12268_15532# sg13g2_nor2b_1_0.Y 0.01673f
C1773 sg13g2_inv_1_1.A a_13936_14726# 0.00238f
C1774 sg13g2_a21oi_1_0.A1 a_13864_16082# 0.00342f
C1775 adc_start sg13g2_dfrbpq_1_1.Q 0.008f
C1776 sg13g2_a21o_1_1.A2 VDD 0.50225f
C1777 sg13g2_a21oi_1_0.A1 a_13679_14845# 0
C1778 a_13866_14020# sg13g2_inv_1_1.Y 0
C1779 uart_busy a_15976_25068# 0.26742f
C1780 a_10024_15996# sg13g2_dfrbpq_1_4.D 0.00179f
C1781 a_14152_5842# sg13g2_buf_1_0.A 0.00233f
C1782 sg13g2_nor2_1_0.B a_12357_13701# 0.00142f
C1783 a_14532_15552# a_15856_16238# 0
C1784 a_14949_15213# a_14859_16007# 0.00237f
C1785 a_16458_14020# sg13g2_inv_1_0.Y 0
C1786 a_14188_17061# sg13g2_inv_1_0.Y 0.01227f
C1787 a_14506_13945# a_14820_13735# 0.00463f
C1788 a_14246_15234# sg13g2_buf_1_0.A 0
C1789 sg13g2_a22oi_1_0.B2 a_15976_25068# 0.24834f
C1790 a_14144_23986# sg13g2_a21oi_1_0.A2 0.00131f
C1791 sg13g2_dfrbpq_1_4.D sg13g2_nor2_1_0.Y 0.22754f
C1792 a_15599_16357# sg13g2_inv_1_1.A 0.00294f
C1793 a_12046_15276# sg13g2_inv_1_0.Y 0.00348f
C1794 sg13g2_buf_1_0.A a_14336_5498# 0.02549f
C1795 sg13g2_inv_1_1.A sg13g2_buf_1_0.A 0.00165f
C1796 sg13g2_a21oi_1_0.A1 a_14235_17564# 0.27988f
C1797 sg13g2_nor2b_1_0.Y a_12297_14113# 0
C1798 sg13g2_a21oi_1_0.A1 a_16266_15996# 0
C1799 a_11654_13722# a_12817_14018# 0
C1800 a_11940_14040# a_12459_13844# 0.34114f
C1801 a_14998_16742# VDD 0.01065f
C1802 a_15791_15311# a_15856_16238# 0
C1803 sg13g2_dfrbpq_1_0.CLK a_12134_14922# 0.00446f
C1804 sg13g2_inv_1_0.Y a_12459_13844# 0.48314f
C1805 sg13g2_dfrbpq_1_5.Q sg13g2_o21ai_1_0.B1 0.00279f
C1806 sg13g2_dfrbpq_1_1.Q a_16051_14746# 0.22317f
C1807 a_14506_13945# sg13g2_and2_1_0.X 0.00937f
C1808 a_12357_13701# a_13456_13942# 0
C1809 a_12459_13844# a_13199_13799# 0.26905f
C1810 a_12537_16119# sg13g2_dfrbpq_1_0.CLK 0
C1811 a_13864_16082# a_13029_16725# 0.00104f
C1812 a_25672_11890# VDD 0.00121f
C1813 a_25856_16668# VDD 0
C1814 sg13g2_dfrbpq_1_0.CLK a_13297_14837# 0.00575f
C1815 a_14757_16007# a_14912_16878# 0.00112f
C1816 a_15217_15998# a_14054_16434# 0
C1817 sg13g2_inv_1_0.Y a_13516_14037# 0.01414f
C1818 a_14155_12256# sg13g2_buf_1_4.A 0.00395f
C1819 sg13g2_dfrbpq_1_3.D a_13936_14726# 0
C1820 a_12326_16746# sg13g2_a21oi_1_0.A2 0.00214f
C1821 a_13199_13799# a_13516_14037# 0.00247f
C1822 a_14859_16007# sg13g2_dfrbpq_1_0.CLK 0.0562f
C1823 sg13g2_dfrbpq_1_0.CLK a_12777_14531# 0
C1824 a_12335_16357# a_12134_14922# 0
C1825 a_14073_17061# sg13g2_a21oi_1_0.A2 0.00165f
C1826 a_13664_10830# VDD 0.06411f
C1827 a_11914_13945# a_11654_13722# 0.75507f
C1828 a_16735_15972# sg13g2_a21o_1_1.A2 0.00131f
C1829 wake_up_sg a_11595_16007# 0
C1830 a_16832_15366# sg13g2_dfrbpq_1_3.Q 0.01342f
C1831 sg13g2_dfrbpq_1_3.D a_15599_16357# 0
C1832 a_14246_13722# a_14346_14484# 0
C1833 sg13g2_dfrbpq_1_3.D sg13g2_buf_1_0.A 0.00454f
C1834 sg13g2_inv_1_0.Y a_9728_13854# 0.00154f
C1835 a_14697_16043# VDD 0
C1836 a_13480_10830# sg13g2_buf_1_4.A 0.00195f
C1837 a_12046_15276# a_12134_14922# 0
C1838 a_12652_16119# a_12592_16238# 0.01042f
C1839 a_12537_16119# a_12335_16357# 0.00689f
C1840 a_13131_16868# sg13g2_dfrbpq_1_4.D 0
C1841 Timer_en a_13960_4782# 0.01683f
C1842 a_14144_23986# VDD 0.00293f
C1843 a_14340_16000# sg13g2_dfrbpq_1_6.D 0.0053f
C1844 sg13g2_dfrbpq_1_3.Q sg13g2_dfrbpq_1_5.Q 0.46867f
C1845 sg13g2_inv_2_1.A a_17696_15156# 0
C1846 a_15409_15530# VDD 0.0077f
C1847 a_14144_17594# sg13g2_inv_1_0.Y 0
C1848 a_14061_12256# a_13838_12256# 0
C1849 a_14340_16000# sg13g2_o21ai_1_0.A1 0.00316f
C1850 a_12652_16119# sg13g2_nor2_1_0.B 0
C1851 sg13g2_nor2_1_0.B a_12939_14495# 0.00444f
C1852 sg13g2_a22oi_1_0.B2 a_14757_16007# 0.04061f
C1853 a_14628_16421# sg13g2_dfrbpq_1_6.D 0.0029f
C1854 a_16458_15532# VDD 0.38282f
C1855 sg13g2_inv_1_0.Y a_12394_14452# 0.27901f
C1856 a_14061_12256# a_14152_10736# 0
C1857 sg13g2_inv_1_1.A a_15784_14570# 0
C1858 wake_up_sg sg13g2_inv_1_0.Y 0.00145f
C1859 a_12357_13701# a_12939_14495# 0
C1860 sg13g2_a21oi_1_0.A1 a_13864_16426# 0.00382f
C1861 sg13g2_dfrbpq_1_4.D a_11595_16007# 0.02579f
C1862 sg13g2_nor2_1_0.B a_13297_14486# 0
C1863 sg13g2_dfrbpq_1_6.D sg13g2_a21oi_1_0.A2 0.05283f
C1864 a_12326_16746# VDD 0.7807f
C1865 sg13g2_a22oi_1_0.B2 a_15217_16349# 0.00677f
C1866 a_16210_15234# VDD 0
C1867 sg13g2_o21ai_1_0.A1 sg13g2_a21oi_1_0.A2 0
C1868 a_11914_13945# sg13g2_a21o_1_0.X 0.00113f
C1869 a_14073_17061# VDD 0.00274f
C1870 sg13g2_inv_1_0.Y a_13936_14726# 0.10353f
C1871 a_15791_15311# a_16051_14746# 0
C1872 a_11940_14040# sg13g2_buf_1_0.A 0.00175f
C1873 a_13866_14020# sg13g2_dfrbpq_1_0.CLK 0.00307f
C1874 a_13199_13799# a_13936_14726# 0
C1875 a_13456_13942# a_12939_14495# 0
C1876 sg13g2_and2_1_0.X a_14346_14484# 0
C1877 sg13g2_dfrbpq_1_4.D a_11953_15998# 0.00363f
C1878 a_15599_16357# sg13g2_inv_1_0.Y 0.13423f
C1879 a_15096_17064# VDD 0.01832f
C1880 sg13g2_inv_1_0.Y sg13g2_buf_1_0.A 0.69243f
C1881 a_13768_10736# a_13664_10620# 0
C1882 a_13480_10830# a_13664_10830# 0.0524f
C1883 a_13199_13799# sg13g2_buf_1_0.A 0.0145f
C1884 adc_start a_15051_13844# 0
C1885 a_15697_15311# sg13g2_a21o_1_1.A2 0
C1886 a_11302_16421# VDD 0
C1887 sg13g2_dfrbpq_1_6.D a_14148_16434# 0
C1888 a_12612_17064# sg13g2_inv_1_1.Y 0
C1889 a_14538_17044# a_14314_15964# 0
C1890 sg13g2_dfrbpq_1_3.D a_15784_14570# 0.02888f
C1891 sg13g2_dfrbpq_1_0.CLK a_15784_14914# 0.00347f
C1892 sg13g2_inv_1_0.Y sg13g2_dfrbpq_1_4.D 0.15656f
C1893 a_13618_13722# VDD 0
C1894 sg13g2_buf_1_6.X a_9728_13854# 0.02132f
C1895 a_14340_16000# sg13g2_o21ai_1_0.B1 0
C1896 clk_gating_en VDD 0.20604f
C1897 a_14440_5412# sc_en 0.24441f
C1898 a_12134_14922# a_12394_14452# 0.75507f
C1899 a_12241_16357# VDD 0
C1900 sg13g2_inv_1_1.A sg13g2_nor2_1_0.Y 0
C1901 sg13g2_a22oi_1_0.B2 a_14314_15964# 0.00142f
C1902 a_13105_13799# a_13618_13722# 0
C1903 adc_done adc_start 0.00514f
C1904 sg13g2_dfrbpq_1_6.D VDD 0.58292f
C1905 a_14532_14040# sg13g2_dfrbpq_1_1.Q 0
C1906 a_14949_13701# a_15784_14570# 0.00171f
C1907 a_15993_14037# VDD 0
C1908 a_14628_16421# sg13g2_o21ai_1_0.B1 0
C1909 a_12268_15532# VDD 0.00713f
C1910 a_14912_16668# sg13g2_dfrbpq_1_0.CLK 0
C1911 sg13g2_o21ai_1_0.A1 VDD 0.45976f
C1912 a_14248_4688# a_13960_4782# 0.00536f
C1913 a_14246_15234# sg13g2_inv_1_1.A 0.02125f
C1914 a_12420_14488# a_12708_14909# 0.43707f
C1915 a_14248_23556# tx_start 0.2541f
C1916 a_14532_15552# sg13g2_a21oi_1_0.A1 0
C1917 adc_start a_15697_13799# 0
C1918 a_15688_25498# VDD 0.00207f
C1919 a_16210_13722# sg13g2_and2_1_0.X 0
C1920 a_14912_16878# a_14998_16742# 0
C1921 sg13g2_o21ai_1_0.B1 sg13g2_a21oi_1_0.A2 0.0284f
C1922 a_14246_15234# a_14340_15234# 0.00716f
C1923 a_15051_15356# a_15409_15530# 0.02138f
C1924 a_14340_16000# a_14566_16421# 0.0052f
C1925 a_15791_13799# sg13g2_dfrbpq_1_1.Q 0.0075f
C1926 a_12228_13735# a_11940_14040# 0.43707f
C1927 a_25856_17938# VDD 0
C1928 a_17024_13644# VDD 0
C1929 a_14506_13945# VDD 0.10142f
C1930 a_7816_15996# sg13g2_dfrbpq_1_0.CLK 0.2561f
C1931 a_12394_14452# a_12777_14531# 0.00333f
C1932 a_12837_14495# a_13585_14845# 0.01058f
C1933 sg13g2_nor2_1_0.A a_12612_17064# 0
C1934 a_12297_14113# VDD 0
C1935 timer_done sg13g2_buf_1_0.A 0.34877f
C1936 a_12228_13735# sg13g2_inv_1_0.Y 0.01622f
C1937 a_17128_13760# sg13g2_a21o_1_1.A2 0
C1938 sg13g2_dfrbpq_1_5.Q a_15680_16668# 0.0013f
C1939 sg13g2_buf_1_0.A a_14632_4688# 0.24846f
C1940 a_12650_15532# sg13g2_nor2_1_0.A 0
C1941 a_13401_14037# a_13456_13942# 0.00412f
C1942 a_13131_16868# sg13g2_nor2_1_0.Y 0.00365f
C1943 a_14246_15234# a_14820_15247# 0.31978f
C1944 a_14340_16000# sg13g2_dfrbpq_1_3.Q 0
C1945 a_14566_16421# a_14628_16421# 0
C1946 sg13g2_a21oi_1_0.A1 a_13871_16823# 0.01324f
C1947 uart_done sg13g2_a21oi_1_0.A2 0.03225f
C1948 a_14820_15247# sg13g2_inv_1_1.A 0.0019f
C1949 sg13g2_inv_2_1.A sg13g2_a21o_1_1.A2 0.23726f
C1950 sg13g2_dfrbpq_1_3.D sg13g2_nor2_1_0.Y 0
C1951 a_13679_14845# a_14098_14922# 0.00174f
C1952 a_12939_14495# a_13297_14486# 0.02138f
C1953 sg13g2_a22oi_1_0.B2 sg13g2_a21o_1_1.A2 0
C1954 a_14758_15247# sg13g2_a21oi_1_0.A1 0
C1955 sg13g2_buf_1_5.X a_13768_10736# 0.00702f
C1956 a_14144_23642# a_13960_25068# 0
C1957 a_14566_16421# sg13g2_a21oi_1_0.A2 0
C1958 a_16840_13644# sg13g2_a21o_1_1.A2 0
C1959 a_15791_15311# a_15993_15549# 0.00689f
C1960 a_14859_16007# a_15599_16357# 0.26905f
C1961 a_14538_17044# a_14998_16742# 0
C1962 sg13g2_inv_1_0.Y a_15784_14570# 0
C1963 a_15217_15998# sg13g2_dfrbpq_1_0.CLK 0.00669f
C1964 sg13g2_inv_1_1.A a_13131_16868# 0
C1965 a_14506_15457# a_14532_15552# 0.36952f
C1966 sg13g2_dfrbpq_1_3.D a_14246_15234# 0.28605f
C1967 a_12537_16119# sg13g2_dfrbpq_1_4.D 0.00153f
C1968 sg13g2_dfrbpq_1_4.D a_13297_14837# 0
C1969 sg13g2_dfrbpq_1_3.D sg13g2_inv_1_1.A 0.49583f
C1970 sg13g2_inv_1_0.Y a_13881_14607# 0.00451f
C1971 a_15505_16357# sg13g2_dfrbpq_1_5.Q 0.00389f
C1972 sg13g2_a22oi_1_0.B2 a_14998_16742# 0.10281f
C1973 sg13g2_a21oi_1_0.A1 a_13777_16823# 0.00351f
C1974 a_13856_25154# sg13g2_a21oi_1_0.A2 0
C1975 a_9728_13644# VDD 0
C1976 a_14889_15625# sg13g2_dfrbpq_1_0.CLK 0
C1977 a_13768_10736# Timer_en 0.24441f
C1978 a_11595_16007# sg13g2_nor2_1_0.Y 0
C1979 a_14340_16000# a_14054_16434# 0.41329f
C1980 a_14949_15213# sg13g2_dfrbpq_1_5.Q 0
C1981 sg13g2_dfrbpq_1_3.D a_14340_15234# 0
C1982 a_14859_16007# sg13g2_dfrbpq_1_4.D 0
C1983 a_12166_13735# sg13g2_a21o_1_0.X 0
C1984 sg13g2_o21ai_1_0.B1 VDD 0.6707f
C1985 a_13029_16725# a_13871_16823# 0.00332f
C1986 a_12612_17064# a_14128_16966# 0.00242f
C1987 a_16832_15156# VDD 0
C1988 a_13702_12532# sg13g2_inv_1_0.Y 0
C1989 a_14336_5842# Timer_en 0
C1990 a_13459_12404# a_13838_12256# 0
C1991 a_15697_15311# a_16210_15234# 0
C1992 a_14628_16421# a_14054_16434# 0.31978f
C1993 sg13g2_nor2b_1_0.Y sg13g2_nor2_1_0.A 0.22641f
C1994 sg13g2_dfrbpq_1_3.D a_14820_15247# 0.00833f
C1995 adc_en a_13960_4782# 0.02118f
C1996 sg13g2_a21oi_1_0.A1 a_12592_16238# 0
C1997 a_14314_15964# a_13679_14845# 0
C1998 a_12837_14495# VDD 0.26539f
C1999 a_13029_16725# a_13489_17042# 0.01483f
C2000 a_12612_17064# sg13g2_dfrbpq_1_0.CLK 0.0952f
C2001 sg13g2_inv_1_1.A a_16048_13942# 0
C2002 a_16832_15366# sg13g2_dfrbpq_1_0.CLK 0
C2003 a_10024_15996# sg13g2_inv_1_0.Y 0
C2004 uart_done VDD 0.20954f
C2005 a_13489_16767# a_13131_16868# 0.00104f
C2006 a_12900_16759# sg13g2_dfrbpq_1_0.CLK 0.00481f
C2007 a_13777_16823# a_13029_16725# 0.01058f
C2008 a_16294_14484# VDD 0.37801f
C2009 a_14054_16434# sg13g2_a21oi_1_0.A2 0.00243f
C2010 a_14144_4782# VDD 0.06713f
C2011 a_13866_14020# a_13936_14726# 0
C2012 a_13105_13799# a_12837_14495# 0
C2013 a_15791_15311# a_15791_13799# 0
C2014 sg13g2_inv_1_0.Y sg13g2_nor2_1_0.Y 0.75458f
C2015 sg13g2_a21oi_1_0.A1 sg13g2_nor2_1_0.B 0
C2016 a_15051_15356# sg13g2_o21ai_1_0.A1 0
C2017 a_14566_16421# VDD 0
C2018 a_12326_16746# a_11493_16007# 0
C2019 a_14346_14484# VDD 0.40857f
C2020 tx_start a_15872_25498# 0
C2021 a_14246_13722# sg13g2_dfrbpq_1_0.CLK 0.00363f
C2022 sg13g2_dfrbpq_1_5.Q sg13g2_dfrbpq_1_0.CLK 0.00304f
C2023 a_15409_15530# sg13g2_a22oi_1_0.B2 0.00156f
C2024 a_14246_15234# sg13g2_inv_1_0.Y 0.11855f
C2025 a_13866_14020# sg13g2_buf_1_0.A 0.05756f
C2026 sg13g2_buf_1_4.A a_13679_14845# 0
C2027 a_13856_25154# VDD 0.09174f
C2028 reset sg13g2_inv_1_0.Y 0
C2029 a_16840_13854# sg13g2_a21o_1_1.A2 0.0012f
C2030 sg13g2_dfrbpq_1_3.Q VDD 0.64661f
C2031 a_14340_16000# sg13g2_inv_1_1.Y 0.00528f
C2032 a_10790_16434# a_11050_15964# 0.75507f
C2033 a_13192_12132# sg13g2_a21o_1_0.X 0.00379f
C2034 sg13g2_dfrbpq_1_3.D a_14949_13701# 0.00226f
C2035 sg13g2_dfrbpq_1_0.CLK a_11364_16421# 0.00868f
C2036 a_12612_17064# a_12335_16357# 0.00248f
C2037 sg13g2_inv_1_1.A sg13g2_inv_1_0.Y 0.07242f
C2038 a_12136_16878# a_12326_16746# 0.00201f
C2039 a_12900_16759# a_12335_16357# 0
C2040 a_16458_15532# sg13g2_inv_2_1.A 0.00627f
C2041 a_16458_15532# sg13g2_a22oi_1_0.B2 0.00158f
C2042 a_14054_16434# a_14148_16434# 0.00716f
C2043 a_14340_15234# sg13g2_inv_1_0.Y 0
C2044 a_14246_13722# a_15409_14018# 0
C2045 a_14532_14040# a_15051_13844# 0.34114f
C2046 a_15697_15311# sg13g2_o21ai_1_0.A1 0
C2047 a_14628_16421# sg13g2_inv_1_1.Y 0
C2048 sg13g2_nor2_1_0.A a_11464_13854# 0
C2049 sg13g2_dfrbpq_1_0.CLK a_12754_16434# 0
C2050 a_11076_16000# a_11364_16421# 0.43707f
C2051 sg13g2_dfrbpq_1_3.D a_16048_13942# 0
C2052 a_13029_16725# sg13g2_nor2_1_0.B 0.00197f
C2053 a_15856_16238# a_16051_14746# 0
C2054 reset a_8776_13854# 0.03394f
C2055 sg13g2_inv_1_0.Y a_12420_16746# 0
C2056 a_14820_13735# sg13g2_dfrbpq_1_0.CLK 0
C2057 a_14506_15457# sg13g2_nor2_1_0.B 0
C2058 uart_done a_13856_25498# 0.00127f
C2059 sg13g2_inv_1_1.Y sg13g2_a21oi_1_0.A2 0.02467f
C2060 a_14912_16878# sg13g2_dfrbpq_1_6.D 0.0023f
C2061 a_14820_15247# sg13g2_inv_1_0.Y 0.00549f
C2062 a_14054_16434# VDD 0.80787f
C2063 sg13g2_nor2b_1_0.Y sg13g2_dfrbpq_1_0.CLK 0
C2064 sg13g2_dfrbpq_1_3.D a_15409_13743# 0
C2065 wake_up_sg a_7816_15996# 0.01128f
C2066 a_11050_15964# a_11433_16043# 0.00333f
C2067 a_14949_13701# a_16048_13942# 0
C2068 a_15051_13844# a_15791_13799# 0.26905f
C2069 a_11493_16007# a_12241_16357# 0.01058f
C2070 sg13g2_o21ai_1_0.A1 a_14912_16878# 0.02686f
C2071 sg13g2_dfrbpq_1_6.D a_11493_16007# 0.00154f
C2072 sg13g2_nor2_1_0.Y a_12134_14922# 0
C2073 a_14859_16007# a_15680_16878# 0.00105f
C2074 a_16210_13722# VDD 0
C2075 sg13g2_inv_1_0.Y a_13131_16868# 0.42194f
C2076 a_13459_12404# sg13g2_dfrbpq_1_0.CLK 0
C2077 a_14061_12256# sg13g2_buf_1_0.A 0
C2078 sg13g2_nor2b_1_0.Y a_11076_16000# 0.00296f
C2079 a_13489_16767# sg13g2_inv_1_0.Y 0
C2080 sg13g2_and2_1_0.X sg13g2_dfrbpq_1_0.CLK 0
C2081 sg13g2_a22oi_1_0.B2 a_15096_17064# 0.01073f
C2082 a_14152_5842# timer_done 0.00274f
C2083 a_12335_16357# a_12754_16434# 0.00174f
C2084 sg13g2_dfrbpq_1_3.Q a_16735_15972# 0.02037f
C2085 sg13g2_dfrbpq_1_3.D sg13g2_inv_1_0.Y 0.12721f
C2086 a_15051_15356# sg13g2_o21ai_1_0.B1 0
C2087 a_11595_16007# a_11953_15998# 0.02138f
C2088 a_15791_13799# a_16108_14037# 0.00247f
C2089 a_14532_14040# a_15697_13799# 0.43239f
C2090 a_14949_13701# a_15409_13743# 0.02396f
C2091 sg13g2_dfrbpq_1_6.D a_13002_15996# 0.00209f
C2092 a_14340_16000# a_15505_16357# 0.43239f
C2093 sg13g2_nor2_1_0.Y a_13297_14837# 0
C2094 timer_done a_14336_5498# 0.00114f
C2095 a_12136_16878# sg13g2_dfrbpq_1_6.D 0.03359f
C2096 a_12817_13743# VDD 0.0013f
C2097 sg13g2_nor2b_1_0.Y a_12335_16357# 0
C2098 a_14949_13701# sg13g2_inv_1_0.Y 0.03758f
C2099 a_14532_15552# a_14757_16007# 0
C2100 a_14949_15213# a_14340_16000# 0
C2101 a_14538_17044# sg13g2_dfrbpq_1_6.D 0.01463f
C2102 a_15791_13799# a_15697_13799# 0.28931f
C2103 a_14506_13945# a_14889_14113# 0.00333f
C2104 a_14152_5498# a_14144_4782# 0
C2105 a_14538_17044# sg13g2_o21ai_1_0.A1 0.00167f
C2106 a_12046_15276# sg13g2_nor2b_1_0.Y 0.30331f
C2107 sg13g2_inv_1_0.Y a_11595_16007# 0.4356f
C2108 reset sg13g2_buf_1_6.X 0.00507f
C2109 sg13g2_a22oi_1_0.B2 sg13g2_dfrbpq_1_6.D 0.10701f
C2110 uart_busy a_15688_25498# 0.00347f
C2111 sg13g2_nor2_1_0.B a_11654_13722# 0
C2112 a_13480_10620# sg13g2_buf_1_0.A 0.00274f
C2113 a_16048_13942# sg13g2_inv_1_0.Y 0.10167f
C2114 sc_en sg13g2_buf_1_0.A 0.17176f
C2115 sg13g2_inv_1_1.Y VDD 0.58576f
C2116 a_17024_13644# a_17128_13760# 0
C2117 sg13g2_a22oi_1_0.B2 sg13g2_o21ai_1_0.A1 0.28907f
C2118 a_14859_16007# sg13g2_inv_1_1.A 0.00517f
C2119 sg13g2_a22oi_1_0.B2 a_15688_25498# 0
C2120 sg13g2_a21oi_1_0.A1 a_15856_16238# 0
C2121 a_11654_13722# a_12357_13701# 0.02454f
C2122 sg13g2_inv_1_0.Y a_11953_15998# 0.01783f
C2123 tx_start sg13g2_a21oi_1_0.A2 0.10845f
C2124 a_15976_25068# a_15872_25154# 0.00624f
C2125 a_14912_16878# sg13g2_o21ai_1_0.B1 0
C2126 a_15916_16119# VDD 0.00728f
C2127 sg13g2_inv_1_0.Y a_11940_14040# 0.41511f
C2128 a_11940_14040# a_13199_13799# 0.01529f
C2129 sg13g2_dfrbpq_1_1.Q sg13g2_a21o_1_1.A2 0.01021f
C2130 a_15680_16668# VDD 0
C2131 a_14340_16000# sg13g2_dfrbpq_1_0.CLK 0.11238f
C2132 a_13838_12256# VDD 0
C2133 a_16108_15549# sg13g2_dfrbpq_1_3.Q 0
C2134 a_16458_15532# a_16266_15996# 0
C2135 sg13g2_inv_1_0.Y a_13199_13799# 0.15132f
C2136 a_14128_16966# sg13g2_a21oi_1_0.A2 0.0045f
C2137 a_14628_16421# sg13g2_dfrbpq_1_0.CLK 0.00448f
C2138 a_12652_16119# a_10790_16434# 0
C2139 a_14152_10736# VDD 0.24333f
C2140 sg13g2_nor2_1_0.A VDD 0.89006f
C2141 a_15697_15311# sg13g2_dfrbpq_1_3.Q 0
C2142 sg13g2_dfrbpq_1_0.CLK a_13585_14845# 0.00879f
C2143 a_14437_17878# sg13g2_dfrbpq_1_6.D 0
C2144 a_13768_10736# sg13g2_buf_1_4.A 0.26372f
C2145 a_14538_17044# sg13g2_o21ai_1_0.B1 0.00196f
C2146 sg13g2_inv_1_0.Y a_8776_13854# 0
C2147 sg13g2_dfrbpq_1_0.CLK sg13g2_a21oi_1_0.A2 0.21854f
C2148 a_15505_16357# VDD 0.00179f
C2149 a_12537_16119# a_11595_16007# 0
C2150 a_25768_25498# VDD 0.00121f
C2151 Timer_en a_13472_4782# 0
C2152 a_14290_16746# sg13g2_a21oi_1_0.A2 0
C2153 a_12612_17064# sg13g2_dfrbpq_1_4.D 0
C2154 a_11914_13945# a_12297_14113# 0.00333f
C2155 sg13g2_a21o_1_0.X a_12357_13701# 0.00165f
C2156 a_14440_5412# VDD 0.26621f
C2157 sg13g2_a22oi_1_0.B2 sg13g2_o21ai_1_0.B1 0.84375f
C2158 sg13g2_inv_1_1.A a_13866_14020# 0
C2159 a_15599_16357# sg13g2_dfrbpq_1_5.Q 0.00807f
C2160 tx_start VDD 0.71931f
C2161 a_14949_15213# VDD 0.25572f
C2162 a_12650_15532# sg13g2_dfrbpq_1_4.D 0
C2163 a_14246_13722# sg13g2_buf_1_0.A 0.03879f
C2164 a_14061_12256# a_13702_12532# 0.01325f
C2165 sg13g2_nor2b_1_0.Y a_12394_14452# 0
C2166 a_13871_16823# a_14314_15964# 0
C2167 sg13g2_a21o_1_0.X a_13456_13942# 0
C2168 sg13g2_nor2_1_0.B a_12708_14909# 0.00303f
C2169 a_13864_16082# sg13g2_dfrbpq_1_6.D 0
C2170 a_16048_15454# VDD 0.16077f
C2171 a_14340_13722# sg13g2_buf_1_0.A 0
C2172 sg13g2_inv_1_0.Y a_12134_14922# 0.1319f
C2173 a_14128_16966# VDD 0.18514f
C2174 sg13g2_dfrbpq_1_4.D a_11364_16421# 0
C2175 a_12537_16119# sg13g2_inv_1_0.Y 0.0058f
C2176 a_14188_17061# sg13g2_a21oi_1_0.A2 0.00197f
C2177 a_14235_17564# sg13g2_dfrbpq_1_6.D 0.00109f
C2178 a_15409_15255# VDD 0.00121f
C2179 sg13g2_inv_1_0.Y a_13297_14837# 0.00217f
C2180 sg13g2_and2_1_0.X a_13936_14726# 0
C2181 a_15791_15311# sg13g2_a21o_1_1.A2 0.00424f
C2182 sg13g2_inv_1_0.Y sg13g2_buf_1_6.X 0.12144f
C2183 sg13g2_dfrbpq_1_3.Q sg13g2_inv_2_1.A 0.11219f
C2184 sg13g2_dfrbpq_1_0.CLK VDD 1.90753f
C2185 sg13g2_a22oi_1_0.B2 sg13g2_dfrbpq_1_3.Q 0.14335f
C2186 a_16458_15532# sg13g2_dfrbpq_1_1.Q 0.00135f
C2187 a_14859_16007# sg13g2_inv_1_0.Y 0.426f
C2188 a_14290_16746# VDD 0.00129f
C2189 sg13g2_inv_1_0.Y a_12777_14531# 0
C2190 a_13768_10736# a_13664_10830# 0.00624f
C2191 a_14437_17878# sg13g2_o21ai_1_0.B1 0.00593f
C2192 a_13459_12404# sg13g2_buf_1_0.A 0.23676f
C2193 a_13105_13799# sg13g2_dfrbpq_1_0.CLK 0.01254f
C2194 sg13g2_nor2b_1_0.Y sg13g2_dfrbpq_1_4.D 0.00483f
C2195 sg13g2_and2_1_0.X sg13g2_buf_1_0.A 0.34242f
C2196 a_11076_16000# VDD 0.07813f
C2197 adc_start a_14532_14040# 0
C2198 sg13g2_buf_1_6.X a_8776_13854# 0
C2199 a_8968_13760# a_8776_13644# 0
C2200 a_15409_14018# VDD 0.00775f
C2201 a_14538_17044# a_14054_16434# 0
C2202 sg13g2_dfrbpq_1_3.D a_15784_14914# 0.00732f
C2203 adc_start a_15791_13799# 0
C2204 a_15505_16357# a_16018_16434# 0
C2205 a_12335_16357# VDD 0.17199f
C2206 sg13g2_a22oi_1_0.B2 a_14054_16434# 0.00267f
C2207 timer_done a_14632_4688# 0.02458f
C2208 a_16458_14020# VDD 0.38571f
C2209 a_14440_5412# a_14152_5498# 0.00524f
C2210 a_13576_4688# a_13472_4572# 0
C2211 a_14188_17061# VDD 0.01393f
C2212 a_12420_14488# a_12837_14495# 0.37583f
C2213 a_12046_15276# VDD 0.21597f
C2214 a_15217_15998# sg13g2_inv_1_1.A 0.00186f
C2215 a_12969_17137# sg13g2_nor2_1_0.Y 0
C2216 a_14949_15213# a_15051_15356# 0.47622f
C2217 a_14144_17594# sg13g2_a21oi_1_0.A2 0.02323f
C2218 a_14532_15552# a_15409_15530# 0
C2219 a_14246_15234# a_14889_15625# 0.00801f
C2220 power_on VSS 0.06665f
C2221 clk_gating_en VSS 1.21618f
C2222 uart_en VSS 0.70739f
C2223 adc_en VSS 1.23599f
C2224 sc_en VSS 0.67035f
C2225 Timer_en VSS 1.20789f
C2226 timer_done VSS 2.12396f
C2227 adc_start VSS 4.4762f
C2228 reset VSS 2.58111f
C2229 adc_done VSS 3.38427f
C2230 wake_up_sg VSS 1.88149f
C2231 clk VSS 2.61586f
C2232 tx_start VSS 1.6554f
C2233 uart_busy VSS 1.76724f
C2234 uart_done VSS 1.51195f
C2235 VDD VSS 1.38739p
C2236 a_25768_4572# VSS 0.02451f $ **FLOATING
C2237 a_25768_4782# VSS 0.1466f $ **FLOATING
C2238 a_14144_4572# VSS 0.00582f $ **FLOATING
C2239 a_13960_4572# VSS 0.01837f $ **FLOATING
C2240 a_14144_4782# VSS 0.03789f $ **FLOATING
C2241 a_13960_4782# VSS 0.08475f $ **FLOATING
C2242 a_13472_4572# VSS 0.00918f $ **FLOATING
C2243 a_13472_4782# VSS 0.06097f $ **FLOATING
C2244 a_14632_4688# VSS 0.36578f
C2245 a_14248_4688# VSS 0.36097f
C2246 a_13576_4688# VSS 0.3804f
C2247 a_14336_5498# VSS 0.03748f $ **FLOATING
C2248 a_14152_5498# VSS 0.09803f $ **FLOATING
C2249 a_14440_5412# VSS 0.37955f
C2250 a_14336_5842# VSS 0.00677f $ **FLOATING
C2251 a_14152_5842# VSS 0.02583f $ **FLOATING
C2252 a_13664_10620# VSS 0.00677f $ **FLOATING
C2253 a_13480_10620# VSS 0.02583f $ **FLOATING
C2254 a_13664_10830# VSS 0.03807f $ **FLOATING
C2255 a_13480_10830# VSS 0.09895f $ **FLOATING
C2256 a_14152_10736# VSS 0.36228f
C2257 a_13768_10736# VSS 0.36904f
C2258 a_25856_11546# VSS 0.07765f $ **FLOATING
C2259 a_25672_11546# VSS 0.09948f $ **FLOATING
C2260 a_25856_11890# VSS 0.00533f $ **FLOATING
C2261 a_25672_11890# VSS 0.02391f $ **FLOATING
C2262 a_14155_12256# VSS 0.00659f
C2263 a_13838_12256# VSS 0.01083f
C2264 a_13192_12132# VSS 0.02473f $ **FLOATING
C2265 a_13702_12532# VSS 0.02782f
C2266 a_13192_12342# VSS 0.09162f $ **FLOATING
C2267 a_14061_12256# VSS 0.30041f
C2268 sg13g2_buf_1_5.X VSS 1.23387f
C2269 sg13g2_a21o_1_0.A2 VSS 0.9063f
C2270 a_13459_12404# VSS 0.51073f
C2271 a_17024_13644# VSS 0.00585f $ **FLOATING
C2272 a_16840_13644# VSS 0.01821f $ **FLOATING
C2273 a_17024_13854# VSS 0.03753f $ **FLOATING
C2274 a_16840_13854# VSS 0.07982f $ **FLOATING
C2275 a_16210_13722# VSS 0.00329f
C2276 a_15697_13799# VSS 0.09498f
C2277 a_15409_13743# VSS 0.00443f
C2278 a_14820_13735# VSS 0.03599f
C2279 a_17128_13760# VSS 0.36807f
C2280 a_16458_14020# VSS 0.41792f
C2281 a_16048_13942# VSS 0.24416f
C2282 a_15791_13799# VSS 0.51893f
C2283 a_14340_13722# VSS 0
C2284 a_13618_13722# VSS 0.00329f
C2285 a_15051_13844# VSS 0.3698f
C2286 a_14949_13701# VSS 0.77467f
C2287 a_14532_14040# VSS 1.57593f
C2288 a_14246_13722# VSS 0.17149f
C2289 sg13g2_and2_1_0.X VSS 0.72237f
C2290 a_14506_13945# VSS 0.23698f
C2291 sg13g2_buf_1_4.A VSS 1.36477f
C2292 a_13105_13799# VSS 0.09495f
C2293 a_12817_13743# VSS 0.00443f
C2294 a_12228_13735# VSS 0.03599f
C2295 a_13866_14020# VSS 0.42028f
C2296 a_13456_13942# VSS 0.24478f
C2297 a_13199_13799# VSS 0.51866f
C2298 a_11748_13722# VSS 0
C2299 a_11464_13644# VSS 0.02444f $ **FLOATING
C2300 a_12459_13844# VSS 0.37091f
C2301 a_12357_13701# VSS 0.77689f
C2302 a_11940_14040# VSS 1.57458f
C2303 a_11654_13722# VSS 0.18412f
C2304 sg13g2_a21o_1_0.X VSS 1.01442f
C2305 a_11464_13854# VSS 0.10225f $ **FLOATING
C2306 a_9728_13644# VSS 0.01015f $ **FLOATING
C2307 a_11914_13945# VSS 0.24067f
C2308 a_9728_13854# VSS 0.04605f $ **FLOATING
C2309 a_8776_13644# VSS 0.02767f $ **FLOATING
C2310 a_8776_13854# VSS 0.10459f $ **FLOATING
C2311 sg13g2_buf_1_6.X VSS 0.70151f
C2312 a_8968_13760# VSS 0.38272f
C2313 a_25768_14570# VSS 0.12848f $ **FLOATING
C2314 a_16294_14484# VSS 0.02632f
C2315 a_25768_14914# VSS 0.02373f $ **FLOATING
C2316 a_16430_14832# VSS 0.01108f
C2317 sg13g2_dfrbpq_1_1.Q VSS 0.79056f
C2318 a_15784_14570# VSS 0.08916f $ **FLOATING
C2319 a_16051_14746# VSS 0.50965f
C2320 a_15784_14914# VSS 0.02464f $ **FLOATING
C2321 sg13g2_buf_1_0.A VSS 3.14746f
C2322 a_14098_14922# VSS 0.00329f
C2323 a_13585_14845# VSS 0.09495f
C2324 a_14346_14484# VSS 0.42699f
C2325 a_13679_14845# VSS 0.52303f
C2326 a_13936_14726# VSS 0.242f
C2327 a_12939_14495# VSS 0.36916f
C2328 a_13297_14837# VSS 0.00443f
C2329 a_12708_14909# VSS 0.03599f
C2330 a_12837_14495# VSS 0.77686f
C2331 a_12420_14488# VSS 1.57543f
C2332 a_12394_14452# VSS 0.23774f
C2333 a_12228_14922# VSS 0
C2334 a_12134_14922# VSS 0.20348f
C2335 a_17696_15156# VSS 0.00892f $ **FLOATING
C2336 a_17696_15366# VSS 0.04724f $ **FLOATING
C2337 a_16832_15156# VSS 0.00765f $ **FLOATING
C2338 sg13g2_a21o_1_1.A2 VSS 1.21093f
C2339 a_16832_15366# VSS 0.04127f $ **FLOATING
C2340 a_16210_15234# VSS 0.00329f
C2341 a_15697_15311# VSS 0.09495f
C2342 a_15409_15255# VSS 0.00443f
C2343 a_14820_15247# VSS 0.03599f
C2344 a_17800_15272# VSS 0.37997f
C2345 a_16458_15532# VSS 0.41936f
C2346 a_16048_15454# VSS 0.2428f
C2347 a_15791_15311# VSS 0.5218f
C2348 a_14340_15234# VSS 0
C2349 a_11848_15156# VSS 0.02614f $ **FLOATING
C2350 a_15051_15356# VSS 0.37179f
C2351 a_14949_15213# VSS 0.78001f
C2352 a_14532_15552# VSS 1.57404f
C2353 a_14246_15234# VSS 0.17239f
C2354 sg13g2_dfrbpq_1_3.D VSS 0.61189f
C2355 a_14506_15457# VSS 0.23687f
C2356 a_12650_15532# VSS 0
C2357 sg13g2_nor2b_1_0.Y VSS 0.54646f
C2358 a_12268_15532# VSS 0
C2359 a_11848_15366# VSS 0.08318f $ **FLOATING
C2360 a_12046_15276# VSS 0.36098f
C2361 a_16735_15972# VSS 0.00152f
C2362 a_17006_16388# VSS 0.00578f
C2363 sg13g2_inv_1_1.A VSS 0.42413f
C2364 a_16018_16434# VSS 0.00329f
C2365 a_15505_16357# VSS 0.09498f
C2366 sg13g2_inv_2_1.A VSS 1.40789f
C2367 sg13g2_dfrbpq_1_3.Q VSS 1.2999f
C2368 a_16266_15996# VSS 0.41808f
C2369 a_15599_16357# VSS 0.52252f
C2370 a_15856_16238# VSS 0.24086f
C2371 a_14859_16007# VSS 0.37055f
C2372 a_15217_16349# VSS 0.00443f
C2373 a_14628_16421# VSS 0.03599f
C2374 a_13864_16082# VSS 0.08174f $ **FLOATING
C2375 a_13499_15996# VSS 0.00632f
C2376 a_14757_16007# VSS 0.78589f
C2377 a_14340_16000# VSS 1.57504f
C2378 a_14314_15964# VSS 0.2373f
C2379 a_14148_16434# VSS 0
C2380 a_14054_16434# VSS 0.18236f
C2381 sg13g2_inv_1_1.Y VSS 0.342f
C2382 a_13864_16426# VSS 0.0234f $ **FLOATING
C2383 a_13601_16344# VSS 0.01118f
C2384 sg13g2_nor2_1_0.Y VSS 0.66093f
C2385 sg13g2_nor2_1_0.B VSS 0.93284f
C2386 a_12754_16434# VSS 0.00329f
C2387 a_12241_16357# VSS 0.09499f
C2388 a_13002_15996# VSS 0.42042f
C2389 a_12335_16357# VSS 0.52459f
C2390 a_12592_16238# VSS 0.23909f
C2391 a_11595_16007# VSS 0.37009f
C2392 a_11953_16349# VSS 0.00443f
C2393 a_11364_16421# VSS 0.03599f
C2394 a_11493_16007# VSS 0.77341f
C2395 a_11076_16000# VSS 1.57798f
C2396 a_11050_15964# VSS 0.23857f
C2397 a_10884_16434# VSS 0
C2398 a_10790_16434# VSS 0.20578f
C2399 sg13g2_dfrbpq_1_4.D VSS 0.3693f
C2400 sg13g2_nor2_1_0.A VSS 1.02565f
C2401 a_9920_16082# VSS 0.04735f $ **FLOATING
C2402 a_10024_15996# VSS 0.37713f
C2403 a_9920_16426# VSS 0.00892f $ **FLOATING
C2404 a_7816_15996# VSS 0.38385f
C2405 a_25856_16668# VSS 0.00748f $ **FLOATING
C2406 a_25856_16878# VSS 0.08592f $ **FLOATING
C2407 a_15680_16668# VSS 0.00697f $ **FLOATING
C2408 a_15496_16668# VSS 0.01913f $ **FLOATING
C2409 a_15680_16878# VSS 0.03558f $ **FLOATING
C2410 a_15496_16878# VSS 0.0819f $ **FLOATING
C2411 a_14912_16668# VSS 0.0054f $ **FLOATING
C2412 a_14998_16742# VSS 0.22026f
C2413 sg13g2_dfrbpq_1_5.Q VSS 1.1949f
C2414 a_14912_16878# VSS 0.0424f $ **FLOATING
C2415 a_14290_16746# VSS 0.00329f
C2416 a_13777_16823# VSS 0.095f
C2417 a_13489_16767# VSS 0.00443f
C2418 a_12900_16759# VSS 0.03599f
C2419 sg13g2_o21ai_1_0.A1 VSS 0.5681f
C2420 a_14538_17044# VSS 0.41947f
C2421 a_14128_16966# VSS 0.2437f
C2422 a_13871_16823# VSS 0.51719f
C2423 a_12420_16746# VSS 0
C2424 a_12136_16668# VSS 0.02444f $ **FLOATING
C2425 sg13g2_dfrbpq_1_0.CLK VSS 3.32437f
C2426 a_13131_16868# VSS 0.37453f
C2427 a_13029_16725# VSS 0.79298f
C2428 a_12612_17064# VSS 1.57631f
C2429 a_12326_16746# VSS 0.18395f
C2430 sg13g2_dfrbpq_1_6.D VSS 0.5976f
C2431 a_12136_16878# VSS 0.1023f $ **FLOATING
C2432 sg13g2_inv_1_0.Y VSS 6.6032f
C2433 a_12586_16969# VSS 0.24067f
C2434 a_25856_17594# VSS 0.08592f $ **FLOATING
C2435 a_25856_17938# VSS 0.00748f $ **FLOATING
C2436 sg13g2_o21ai_1_0.B1 VSS 0.57643f
C2437 a_14437_17878# VSS 0.00852f
C2438 a_14144_17594# VSS 0.05786f $ **FLOATING
C2439 a_14235_17564# VSS 0.38895f
C2440 a_14144_17938# VSS 0.00899f $ **FLOATING
C2441 a_25768_23642# VSS 0.12888f $ **FLOATING
C2442 a_25768_23986# VSS 0.02422f $ **FLOATING
C2443 a_14144_23642# VSS 0.06023f $ **FLOATING
C2444 sg13g2_a21oi_1_0.A1 VSS 2.2072f
C2445 a_14248_23556# VSS 0.38693f
C2446 a_14144_23986# VSS 0.00902f $ **FLOATING
C2447 a_25768_25154# VSS 0.14597f $ **FLOATING
C2448 a_25768_25498# VSS 0.02451f $ **FLOATING
C2449 sg13g2_a22oi_1_0.B2 VSS 3.0457f
C2450 a_15872_25154# VSS 0.03985f $ **FLOATING
C2451 a_15688_25154# VSS 0.10206f $ **FLOATING
C2452 a_15976_25068# VSS 0.384f
C2453 a_15872_25498# VSS 0.00693f $ **FLOATING
C2454 a_15688_25498# VSS 0.02637f $ **FLOATING
C2455 sg13g2_a21oi_1_0.A2 VSS 2.71f
C2456 a_13856_25154# VSS 0.04901f $ **FLOATING
C2457 a_13960_25068# VSS 0.38011f
C2458 a_13856_25498# VSS 0.00907f $ **FLOATING
.ends

