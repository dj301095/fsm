* NGSPICE file created from fsm_flat.ext - technology: ihp-sg13

.subckt fsm_flat Timer_en adc_en clk_gating_en power_on sc_en timer_done tx_start
+ uart_busy uart_done uart_en adc_done adc_start clk reset wake_up_sg VDD VSS
X0 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=2.28077n ps=0.01084 w=0.42u l=1u
x1 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=3.17827n ps=0.01242 w=1u l=1u
x2 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x4 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x5 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x6 VSS a_16048_15454# a_15697_15311# VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
x7 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x8 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x9 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x10 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1 u l=1u
x11 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x12 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x13 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x14 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x15 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x16 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x17 a_14697_16043# a_14340_16000# VDD VDD sg13_lv_pmos ad=63f pd=0.72u as=0.1563p ps=1.22u w=0.42u l=0.13u
x18 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x19 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x20 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x21 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x22 a_14054_16434# sg13_inv_1_1.Y VDD VDD sg13_lv_pmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
x23 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x24 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x25 a_11654_13722# a_12459_13844# a_11914_13945# VDD sg13_lv_pmos ad=0.1428p pd=1.52u as=79.8f ps=0.8u w=0.42u l=0.13u
x26 VSS sg13_a21oi_1_0.A1 a_14248_23556# VSS sg13_lv_nmos ad=0.14875p pd=1.16u as=0.187p ps=1.78u w=0.55u l=0.13u
x27 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x28 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x29 VDD sg13_inv_1_0.Y a_12394_14452# VDD sg13_lv_pmos ad=0.1563p pd=1.22u as=0.147p ps=1.54u w=0.42u l=0.13u
x30 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x31 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x32 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x33 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x34 a_16048_13942# sg13_inv_1_0.Y a_16108_14037# VDD sg13_lv_pmos ad=79.8f pd=0.8u as=0.204p ps=1.835u w=0.42u l=0.13u
x35 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x36 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x37 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x38 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x39 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x40 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x41 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x42 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x43 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x44 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x45 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x46 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x47 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x48 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x49 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x50 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x51 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x52 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x53 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x54 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x55 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x56 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x57 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x58 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x59 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x60 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x61 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x62 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x63 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x64 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x65 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x66 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x67 a_13297_14486# a_12837_14495# a_12939_14495# VDD sg13_lv_pmos ad=0.41165p pd=2.12u as=0.3864p ps=2.93u w=1.12u l=0.13u
x68 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x69 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x70 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x71 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x72 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x73 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x74 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x75 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x76 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x77 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x78 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x79 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x80 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x81 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x82 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x83 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x84 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x85 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x86 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x87 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x88 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x89 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x90 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x91 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x92 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x93 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x94 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x95 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x96 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x97 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x98 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x99 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x100 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x101 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x102 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x103 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x104 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x105 sg13_inv_2_1.A a_17800_15272# VDD VDD sg13_lv_pmos ad=0.42p pd=2.99u as=0.2114p ps=1.54u w=1.12u l=0.13u
x106 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x107 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x108 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x109 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x110 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x111 a_14340_13722# sg13_and2_1_0.X a_14246_13722# VSS sg13_lv_nmos ad=60.89999f pd=0.71u as=0.1428p ps=1.52u w=0.42u l=0.13u
x112 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x113 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x114 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x115 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x116 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x117 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x118 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x119 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x120 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x121 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x122 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x123 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x124 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x125 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x126 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x127 a_15217_16349# a_14757_16007# a_14859_16007# VSS sg13_lv_nmos ad=0.31732p pd=1.805u as=0.2516p ps=2.16u w=0.74u l=0.13u
x128 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x129 VSS adc_done a_17800_15272# VSS sg13_lv_nmos ad=0.14875p pd=1.16u as=0.187p ps=1.78u w=0.55u l=0.13u
x130 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x131 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x132 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x133 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x134 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x135 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x136 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x137 a_12708_14909# a_12420_14488# a_12646_14909# VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=37.8f ps=0.6u w=0.42u l=0.13u
x138 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x139 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x140 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x141 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x142 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x143 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x144 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x145 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x146 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x147 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x148 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x149 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x150 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x151 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x152 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x153 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x154 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x155 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x156 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x157 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x158 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x159 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x160 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x161 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x162 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x163 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x164 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x165 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x166 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x167 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x168 a_14340_16000# a_14314_15964# VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0.36237p ps=2.605u w=1u l=0.13u
x169 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x170 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x171 sg13_buf_1_5.X a_14152_10736# VSS VSS sg13_lv_nmos ad=0.2886p pd=2.26u as=0.14875p ps=1.16u w=0.74u l=0.13u
x172 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x173 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x174 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x175 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x176 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x177 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x178 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x179 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x180 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x181 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x182 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x183 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x184 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x185 sg13_a21oi_1_0.A1 a_14538_17044# VSS VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.1406p ps=1.12u w=0.74u l=0.13u
x186 sg13_inv_1_1.A sg13_a22oi_1_0.B2 a_16735_16388# VSS sg13_lv_nmos ad=0.2664p pd=1.46u as=0.13875p ps=1.115u w=0.74u l=0.13u
x187 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x188 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x189 sg13_dfrbpq_1_0.CLK a_7816_15996# VDD VDD sg13_lv_pmos ad=0.42p pd=2.99u as=0.2114p ps=1.54u w=1.12u l=0.13u
x190 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x191 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x192 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x193 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x194 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x195 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x196 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x197 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x198 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x199 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x200 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x201 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x202 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x203 a_13936_14726# sg13_inv_1_0.Y a_13996_14607# VDD sg13_lv_pmos ad=79.8f pd=0.8u as=0.204p ps=1.835u w=0.42u l=0.13u
x204 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x205 a_14314_15964# a_14757_16007# a_14054_16434# VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0.1296p ps=1.52u w=0.42u l=0.13u
x206 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x207 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x208 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x209 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x210 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x211 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x212 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x213 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x214 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x215 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x216 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x217 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x218 sg13_dfrbpq_1_5.Q a_16266_15996# VDD VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
x219 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x220 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x221 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x222 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x223 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x224 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x225 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x226 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x227 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x228 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x229 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x230 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x231 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x232 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x233 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x234 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x235 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x236 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x237 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x238 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x239 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x240 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x241 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x242 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x243 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x244 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x245 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x246 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x247 a_13456_13942# sg13_inv_1_0.Y a_13516_14037# VDD sg13_lv_pmos ad=79.8f pd=0.8u as=0.204p ps=1.835u w=0.42u l=0.13u
x248 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x249 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x250 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x251 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x252 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x253 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x254 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x255 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x256 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x257 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x258 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x259 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x260 VSS sg13_nor2_1_0.B sg13_nor2_1_0.Y VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.1406p ps=1.12u w=0.74u l=0.13u
x261 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x262 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x263 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x264 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x265 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x266 a_13936_14726# a_13679_14845# a_14098_14922# VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=37.8f ps=0.6u w=0.42u l=0.13u
x267 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x268 a_14188_17061# a_14128_16966# a_14073_17061# VDD sg13_lv_pmos ad=0.204p pd=1.835u as=93.45f ps=0.865u w=0.42u l=0.13u
x269 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x270 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x271 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x272 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x273 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x274 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x275 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x276 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x277 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x278 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x279 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x280 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x281 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x282 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x283 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x284 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x285 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x286 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x287 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x288 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x289 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x290 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x291 a_14628_16421# a_14340_16000# a_14566_16421# VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=37.8f ps=0.6u w=0.42u l=0.13u
x292 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x293 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x294 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x295 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x296 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x297 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x298 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x299 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x300 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x301 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x302 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x303 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x304 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x305 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x306 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x307 adc_start a_17128_13760# VDD VDD sg13_lv_pmos ad=0.42p pd=2.99u as=0.2114p ps=1.54u w=1.12u l=0.13u
x308 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x309 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x310 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x311 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x312 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x313 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x314 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x315 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x316 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x317 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x318 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x319 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x320 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x321 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x322 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x323 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x324 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x325 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x326 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x327 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x328 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x329 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x330 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x331 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x332 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x333 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x334 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x335 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x336 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x337 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x338 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x339 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x340 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x341 a_11748_13722# sg13_a21o_1_0.X a_11654_13722# VSS sg13_lv_nmos ad=60.89999f pd=0.71u as=0.1428p ps=1.52u w=0.42u l=0.13u
x342 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x343 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x344 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x345 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x346 a_12612_17064# a_12586_16969# VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0.36237p ps=2.605u w=1u l=0.13u
x347 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x348 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x349 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x350 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x351 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x352 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x353 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x354 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x355 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x356 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x357 a_12646_14909# sg13_inv_1_0.Y VSS VSS sg13_lv_nmos ad=37.8f pd=0.6u as=0.1701p ps=1.65u w=0.42u l=0.13u
x358 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x359 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x360 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x361 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x362 a_12297_14113# a_11940_14040# VDD VDD sg13_lv_pmos ad=63f pd=0.72u as=0.1563p ps=1.22u w=0.42u l=0.13u
x363 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x364 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x365 a_13702_12532# sg13_buf_1_0.A a_13459_12404# VDD sg13_lv_pmos ad=0.2125p pd=1.425u as=0.35p ps=2.7u w=1u l=0.13u
x366 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x367 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x368 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x369 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x370 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x371 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x372 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x373 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x374 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x375 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x376 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x377 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x378 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x379 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x380 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x381 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x382 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x383 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x384 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x385 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x386 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x387 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x388 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x389 a_15409_14018# a_14949_13701# a_15051_13844# VDD sg13_lv_pmos ad=0.41165p pd=2.12u as=0.3864p ps=2.93u w=1.12u l=0.13u
x390 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x391 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x392 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x393 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x394 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x395 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x396 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x397 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x398 adc_en a_13576_4688# VSS VSS sg13_lv_nmos ad=0.2886p pd=2.26u as=0.14875p ps=1.16u w=0.74u l=0.13u
x399 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x400 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x401 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x402 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x403 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x404 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x405 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x406 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x407 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x408 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x409 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x410 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x411 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x412 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x413 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x414 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x415 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x416 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x417 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x418 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x419 VDD reset a_8968_13760# VDD sg13_lv_pmos ad=0.2114p pd=1.54u as=0.2856p ps=2.36u w=0.84u l=0.13u
x420 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x421 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x422 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x423 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x424 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x425 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x426 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x427 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x428 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x429 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x430 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x431 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x432 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x433 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x434 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x435 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x436 VDD a_15791_15311# a_16048_15454# VDD sg13_lv_pmos ad=0.4659p pd=3.65u as=79.8f ps=0.8u w=0.42u l=0.13u
x437 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x438 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x439 VSS a_15599_16357# a_16266_15996# VSS sg13_lv_nmos ad=0.1406p pd=1.12u as=0.2516p ps=2.16u w=0.74u l=0.13u
x440 sg13_inv_1_0.Y sg13_buf_1_6.X VSS VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.2516p ps=2.16u w=0.74u l=0.13u
x441 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x442 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x443 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x444 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x445 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x446 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x447 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x448 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x449 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x450 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x451 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x452 clk_gating_en a_14632_4688# VDD VDD sg13_lv_pmos ad=0.42p pd=2.99u as=0.2114p ps=1.54u w=1.12u l=0.13u
x453 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x454 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x455 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x456 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x457 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x458 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x459 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x460 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x461 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x462 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x463 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x464 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x465 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x466 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x467 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x468 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x469 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x470 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x471 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x472 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x473 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x474 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x475 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x476 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x477 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x478 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x479 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x480 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x481 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x482 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x483 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x484 a_11493_16007# sg13_dfrbpq_1_0.CLK a_11953_16349# VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.31732p ps=1.805u w=0.74u l=0.13u
x485 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x486 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x487 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x488 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x489 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x490 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x491 a_12420_14488# a_12394_14452# VSS VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.1626p ps=1.415u w=0.74u l=0.13u
x492 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x493 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x494 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x495 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x496 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x497 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x498 uart_en a_14248_4688# VSS VSS sg13_lv_nmos ad=0.2886p pd=2.26u as=0.14875p ps=1.16u w=0.74u l=0.13u
x499 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x500 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x501 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x502 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x503 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x504 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x505 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x506 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x507 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x508 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x509 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x510 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x511 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x512 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x513 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x514 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x515 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x516 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x517 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x518 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x519 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x520 a_14340_16000# a_14859_16007# a_15599_16357# VSS sg13_lv_nmos ad=0.3473p pd=2.71u as=0.12665p ps=1.145u w=0.74u l=0.13u
x521 VDD a_15791_13799# a_16458_14020# VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.3864p ps=2.93u w=1.12u l=0.13u
x522 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x523 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x524 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x525 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x526 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x527 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x528 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x529 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x530 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x531 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x532 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x533 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x534 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x535 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x536 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x537 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x538 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x539 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x540 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x541 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x542 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x543 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x544 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x545 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x546 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x547 a_14532_15552# a_14506_15457# VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0.36237p ps=2.605u w=1u l=0.13u
x548 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x549 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x550 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x551 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x552 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x553 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x554 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x555 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x556 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x557 a_14889_14113# a_14532_14040# VDD VDD sg13_lv_pmos ad=63f pd=0.72u as=0.1563p ps=1.22u w=0.42u l=0.13u
x558 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x559 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x560 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x561 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x562 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x563 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x564 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x565 VSS a_12592_16238# a_12241_16357# VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
x566 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x567 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x568 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x569 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x570 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x571 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x572 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x573 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x574 a_14073_17061# a_13131_16868# a_13871_16823# VDD sg13_lv_pmos ad=93.45f pd=0.865u as=0.2048p ps=1.63u w=0.42u l=0.13u
x575 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x576 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x577 a_12586_16969# a_13029_16725# a_12326_16746# VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0.1296p ps=1.52u w=0.42u l=0.13u
x578 a_12592_16238# a_12335_16357# a_12754_16434# VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=37.8f ps=0.6u w=0.42u l=0.13u
x579 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x580 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x581 VSS a_16048_13942# a_15697_13799# VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
x582 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x583 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x584 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x585 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x586 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x587 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x588 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x589 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x590 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x591 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x592 a_11433_16043# a_11076_16000# VDD VDD sg13_lv_pmos ad=63f pd=0.72u as=0.1563p ps=1.22u w=0.42u l=0.13u
x593 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x594 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x595 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x596 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x597 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x598 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x599 a_12817_14018# a_12357_13701# a_12459_13844# VDD sg13_lv_pmos ad=0.41165p pd=2.12u as=0.3864p ps=2.93u w=1.12u l=0.13u
x600 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x601 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x602 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x603 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x604 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x605 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x606 a_14532_15552# a_14506_15457# VSS VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.1626p ps=1.415u w=0.74u l=0.13u
x607 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x608 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x609 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x610 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x611 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x612 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x613 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x614 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x615 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x616 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x617 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x618 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x619 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x620 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x621 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x622 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x623 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x624 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x625 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x626 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x627 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x628 a_13679_14845# a_12837_14495# a_13585_14845# VSS sg13_lv_nmos ad=0.12665p pd=1.145u as=0.1428p ps=1.52u w=0.42u l=0.13u
x629 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x630 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x631 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x632 a_11050_15964# a_11493_16007# a_11433_16043# VDD sg13_lv_pmos ad=79.8f pd=0.8u as=63f ps=0.72u w=0.42u l=0.13u
x633 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x634 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x635 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x636 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x637 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x638 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x639 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x640 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x641 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x642 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x643 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x644 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x645 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x646 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x647 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x648 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x649 a_16735_15972# sg13_dfrbpq_1_3.Q VDD VDD sg13_lv_pmos ad=0.2716p pd=1.605u as=0.3808p ps=2.92u w=1.12u l=0.13u
x650 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x651 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x652 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x653 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x654 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x655 sg13_and2_1_0.X a_14061_12256# VDD VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.1918p ps=1.5u w=1.12u l=0.13u
x656 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x657 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x658 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x659 a_15409_15255# a_14949_15213# a_15051_15356# VSS sg13_lv_nmos ad=0.31732p pd=1.805u as=0.2516p ps=2.16u w=0.74u l=0.13u
x660 a_16051_14746# sg13_dfrbpq_1_1.Q VSS VSS sg13_lv_nmos ad=0.1216p pd=1.02u as=0.15745p ps=1.175u w=0.64u l=0.13u
x661 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x662 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x663 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x664 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x665 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x666 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x667 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x668 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x669 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x670 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x671 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x672 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x673 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x674 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x675 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x676 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x677 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x678 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x679 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x680 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x681 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x682 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x683 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x684 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x685 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x686 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x687 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x688 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x689 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x690 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x691 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x692 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x693 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x694 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x695 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x696 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x697 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x698 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x699 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x700 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x701 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x702 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x703 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x704 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x705 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x706 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x707 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x708 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x709 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x710 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x711 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x712 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x713 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x714 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x715 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x716 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x717 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x718 a_15409_15530# a_14949_15213# a_15051_15356# VDD sg13_lv_pmos ad=0.41165p pd=2.12u as=0.3864p ps=2.93u w=1.12u l=0.13u
x719 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x720 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x721 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x722 VDD a_13199_13799# a_13866_14020# VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.3864p ps=2.93u w=1.12u l=0.13u
x723 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x724 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x725 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x726 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x727 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x728 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x729 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x730 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x731 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x732 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x733 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x734 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x735 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x736 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x737 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x738 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x739 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x740 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x741 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x742 sg13_o21ai_1_0.B1 a_14235_17564# a_14437_17878# VSS sg13_lv_nmos ad=0.333p pd=2.38u as=0.1406p ps=1.12u w=0.74u l=0.13u
x743 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x744 a_12394_14452# a_12837_14495# a_12777_14531# VDD sg13_lv_pmos ad=79.8f pd=0.8u as=63f ps=0.72u w=0.42u l=0.13u
x745 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x746 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x747 VDD sg13_inv_1_0.Y a_14246_13722# VDD sg13_lv_pmos ad=0.36237p pd=2.605u as=79.8f ps=0.8u w=0.42u l=0.13u
x748 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x749 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x750 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x751 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x752 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x753 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x754 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x755 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x756 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x757 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x758 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x759 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x760 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x761 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x762 sc_en a_14440_5412# VSS VSS sg13_lv_nmos ad=0.2886p pd=2.26u as=0.14875p ps=1.16u w=0.74u l=0.13u
x763 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x764 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x765 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x766 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x767 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x768 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x769 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x770 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x771 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x772 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x773 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x774 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x775 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x776 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x777 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x778 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x779 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x780 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x781 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x782 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x783 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x784 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x785 a_13838_12256# sg13_buf_1_4.A a_13459_12404# VSS sg13_lv_nmos ad=81.6f pd=0.895u as=0.1216p ps=1.02u w=0.64u l=0.13u
x786 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x787 VDD a_13871_16823# a_14538_17044# VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.3864p ps=2.93u w=1.12u l=0.13u
x788 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x789 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x790 VSS sg13_inv_1_0.Y a_12228_14922# VSS sg13_lv_nmos ad=0.1626p pd=1.415u as=60.89999f ps=0.71u w=0.42u l=0.13u
x791 VSS a_13456_13942# a_13105_13799# VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
x792 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x793 a_12900_16759# a_13131_16868# a_12586_16969# VSS sg13_lv_nmos ad=0.2373p pd=1.97u as=79.8f ps=0.8u w=0.42u l=0.13u
x794 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x795 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x796 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x797 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x798 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x799 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x800 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x801 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x802 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x803 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x804 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x805 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x806 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x807 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x808 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x809 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x810 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x811 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x812 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x813 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x814 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x815 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x816 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x817 a_14820_15247# a_15051_15356# a_14506_15457# VSS sg13_lv_nmos ad=0.2373p pd=1.97u as=79.8f ps=0.8u w=0.42u l=0.13u
x818 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x819 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x820 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x821 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x822 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x823 sg13_o21ai_1_0.A1 sg13_dfrbpq_1_5.Q VDD VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.3808p ps=2.92u w=1.12u l=0.13u
x824 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x825 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x826 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x827 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x828 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x829 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x830 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x831 a_12969_17137# a_12612_17064# VDD VDD sg13_lv_pmos ad=63f pd=0.72u as=0.1563p ps=1.22u w=0.42u l=0.13u
x832 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x833 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x834 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x835 VSS reset a_8968_13760# VSS sg13_lv_nmos ad=0.14875p pd=1.16u as=0.187p ps=1.78u w=0.55u l=0.13u
x836 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x837 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x838 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x839 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x840 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x841 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x842 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x843 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x844 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x845 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x846 adc_en a_13576_4688# VDD VDD sg13_lv_pmos ad=0.42p pd=2.99u as=0.2114p ps=1.54u w=1.12u l=0.13u
x847 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x848 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x849 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x850 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x851 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x852 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x853 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x854 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x855 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x856 VSS timer_done a_14152_10736# VSS sg13_lv_nmos ad=0.14875p pd=1.16u as=0.187p ps=1.78u w=0.55u l=0.13u
x857 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x858 VSS a_14128_16966# a_13777_16823# VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
x859 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x860 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x861 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x862 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x863 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x864 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x865 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x866 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x867 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x868 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x869 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x870 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x871 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x872 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x873 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x874 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x875 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x876 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x877 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x878 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x879 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x880 sg13_nor2b_1_0.Y a_12046_15276# VSS VSS sg13_lv_nmos ad=0.1406p pd=1.12u as=0.17255p ps=1.25u w=0.74u l=0.13u
x881 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x882 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x883 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x884 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x885 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x886 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x887 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x888 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x889 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x890 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x891 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x892 sg13_dfrbpq_1_3.Q a_16458_15532# VDD VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
x893 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x894 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x895 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x896 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x897 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x898 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x899 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x900 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x901 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x902 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x903 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x904 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x905 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x906 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x907 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x908 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x909 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x910 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x911 a_12420_14488# a_12394_14452# VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0.36237p ps=2.605u w=1u l=0.13u
x912 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x913 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x914 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x915 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x916 a_12537_16119# a_11595_16007# a_12335_16357# VDD sg13_lv_pmos ad=93.45f pd=0.865u as=0.2048p ps=1.63u w=0.42u l=0.13u
x917 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x918 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x919 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x920 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x921 sg13_inv_1_0.Y sg13_buf_1_6.X VDD VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.3808p ps=2.92u w=1.12u l=0.13u
x922 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x923 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x924 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x925 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x926 a_14532_15552# a_15051_15356# a_15791_15311# VSS sg13_lv_nmos ad=0.3473p pd=2.71u as=0.12665p ps=1.145u w=0.74u l=0.13u
x927 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x928 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x929 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x930 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x931 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x932 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x933 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x934 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x935 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x936 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x937 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x938 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x939 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x940 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x941 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x942 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x943 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x944 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x945 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x946 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x947 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x948 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x949 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x950 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x951 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x952 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x953 uart_en a_14248_4688# VDD VDD sg13_lv_pmos ad=0.42p pd=2.99u as=0.2114p ps=1.54u w=1.12u l=0.13u
x954 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x955 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x956 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x957 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x958 sg13_a21o_1_0.A2 sg13_buf_1_5.X VSS VSS sg13_lv_nmos ad=0.1406p pd=1.12u as=0.2516p ps=2.16u w=0.74u l=0.13u
x959 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x960 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x961 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x962 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x963 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x964 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x965 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x966 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x967 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x968 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x969 VDD sg13_inv_1_0.Y a_11654_13722# VDD sg13_lv_pmos ad=0.36237p pd=2.605u as=79.8f ps=0.8u w=0.42u l=0.13u
x970 a_17006_16388# sg13_dfrbpq_1_3.Q sg13_inv_1_1.A VSS sg13_lv_nmos ad=96.2f pd=1u as=0.2664p ps=1.46u w=0.74u l=0.13u
x971 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x972 a_15791_15311# a_14949_15213# a_15697_15311# VSS sg13_lv_nmos ad=0.12665p pd=1.145u as=0.1428p ps=1.52u w=0.42u l=0.13u
x973 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x974 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x975 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x976 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x977 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x978 a_15916_16119# a_15856_16238# a_15801_16119# VDD sg13_lv_pmos ad=0.204p pd=1.835u as=93.45f ps=0.865u w=0.42u l=0.13u
x979 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x980 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x981 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x982 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x983 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x984 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x985 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x986 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x987 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x988 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x989 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x990 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x991 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x992 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x993 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x994 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x995 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x996 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x997 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x998 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x999 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1000 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1001 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1002 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1003 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1004 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1005 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1006 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1007 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1008 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1009 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1010 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1011 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1012 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1013 VDD sg13_buf_1_0.A a_14632_4688# VDD sg13_lv_pmos ad=0.2114p pd=1.54u as=0.2856p ps=2.36u w=0.84u l=0.13u
x1014 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1015 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1016 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1017 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1018 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1019 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1020 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1021 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1022 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1023 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1024 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1025 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1026 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1027 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1028 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1029 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1030 sg13_buf_1_6.X a_8968_13760# VDD VDD sg13_lv_pmos ad=0.42p pd=2.99u as=0.2114p ps=1.54u w=1.12u l=0.13u
x1031 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1032 a_14506_15457# a_14949_15213# a_14246_15234# VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0.1296p ps=1.52u w=0.42u l=0.13u
x1033 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1034 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1035 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1036 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1037 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1038 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1039 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1040 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1041 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1042 a_14820_15247# a_14532_15552# a_14758_15247# VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=37.8f ps=0.6u w=0.42u l=0.13u
x1043 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1044 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1045 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1046 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1047 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1048 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1049 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1050 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1051 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1052 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1053 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1054 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1055 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1056 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1057 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1058 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1059 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1060 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1061 VSS uart_done a_13960_25068# VSS sg13_lv_nmos ad=0.14875p pd=1.16u as=0.187p ps=1.78u w=0.55u l=0.13u
x1062 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1063 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1064 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1065 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1066 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1067 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1068 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1069 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1070 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1071 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1072 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1073 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1074 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1075 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1076 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1077 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1078 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1079 VSS sg13_inv_1_0.Y a_11748_13722# VSS sg13_lv_nmos ad=0.1626p pd=1.415u as=60.89999f ps=0.71u w=0.42u l=0.13u
x1080 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1081 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1082 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1083 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1084 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1085 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1086 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1087 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1088 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1089 a_11076_16000# a_11595_16007# a_12335_16357# VSS sg13_lv_nmos ad=0.3473p pd=2.71u as=0.12665p ps=1.145u w=0.74u l=0.13u
x1090 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1091 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1092 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1093 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1094 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1095 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1096 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1097 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1098 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1099 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1100 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1101 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1102 a_12837_14495# sg13_dfrbpq_1_0.CLK a_13297_14486# VDD sg13_lv_pmos ad=0.4088p pd=2.97u as=0.41165p ps=2.12u w=1.12u l=0.13u
x1103 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1104 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1105 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1106 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1107 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1108 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1109 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1110 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1111 VDD sg13_inv_1_0.Y a_12586_16969# VDD sg13_lv_pmos ad=0.1563p pd=1.22u as=0.147p ps=1.54u w=0.42u l=0.13u
x1112 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1113 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1114 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1115 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1116 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1117 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1118 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1119 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1120 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1121 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1122 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1123 sg13_a22oi_1_0.B2 a_15976_25068# VDD VDD sg13_lv_pmos ad=0.42p pd=2.99u as=0.2114p ps=1.54u w=1.12u l=0.13u
x1124 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1125 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1126 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1127 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1128 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1129 VDD a_14235_17564# sg13_o21ai_1_0.B1 VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
x1130 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1131 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1132 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1133 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1134 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1135 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1136 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1137 a_11953_16349# a_11493_16007# a_11595_16007# VSS sg13_lv_nmos ad=0.31732p pd=1.805u as=0.2516p ps=2.16u w=0.74u l=0.13u
x1138 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1139 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1140 a_12268_15532# a_12046_15276# VDD VDD sg13_lv_pmos ad=0.1176p pd=1.33u as=0.2618p ps=1.63u w=1.12u l=0.13u
x1141 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1142 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1143 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1144 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1145 a_13199_13799# a_12357_13701# a_13105_13799# VSS sg13_lv_nmos ad=0.12665p pd=1.145u as=0.1428p ps=1.52u w=0.42u l=0.13u
x1146 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1147 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1148 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1149 a_13601_16344# sg13_a21oi_1_0.A1 sg13_dfrbpq_1_4.D VSS sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
x1150 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1151 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1152 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1153 a_16018_16434# sg13_inv_1_0.Y VSS VSS sg13_lv_nmos ad=37.8f pd=0.6u as=79.8f ps=0.8u w=0.42u l=0.13u
x1154 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1155 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1156 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1157 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1158 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1159 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1160 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1161 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1162 a_14757_16007# sg13_dfrbpq_1_0.CLK a_15217_16349# VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.31732p ps=1.805u w=0.74u l=0.13u
x1163 a_16210_15234# sg13_inv_1_0.Y VSS VSS sg13_lv_nmos ad=37.8f pd=0.6u as=79.8f ps=0.8u w=0.42u l=0.13u
x1164 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1165 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1166 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1167 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1168 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1169 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1170 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1171 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1172 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1173 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1174 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1175 VDD a_12335_16357# a_13002_15996# VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.3864p ps=2.93u w=1.12u l=0.13u
x1176 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1177 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1178 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1179 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1180 VDD sg13_inv_1_0.Y a_14054_16434# VDD sg13_lv_pmos ad=0.36237p pd=2.605u as=79.8f ps=0.8u w=0.42u l=0.13u
x1181 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1182 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1183 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1184 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1185 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1186 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1187 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1188 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1189 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1190 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1191 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1192 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1193 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1194 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1195 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1196 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1197 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1198 a_14532_14040# a_14506_13945# VSS VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.1626p ps=1.415u w=0.74u l=0.13u
x1199 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1200 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1201 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1202 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1203 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1204 VSS a_16051_14746# sg13_dfrbpq_1_3.D VSS sg13_lv_nmos ad=0.15745p pd=1.175u as=0.2351p ps=2.16u w=0.74u l=0.13u
x1205 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1206 VDD a_15791_13799# a_16048_13942# VDD sg13_lv_pmos ad=0.4659p pd=3.65u as=79.8f ps=0.8u w=0.42u l=0.13u
x1207 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1208 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1209 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1210 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1211 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1212 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1213 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1214 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1215 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1216 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1217 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1218 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1219 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1220 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1221 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1222 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1223 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1224 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1225 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1226 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1227 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1228 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1229 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1230 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1231 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1232 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1233 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1234 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1235 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1236 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1237 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1238 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1239 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1240 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1241 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1242 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1243 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1244 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1245 VSS sg13_buf_1_0.A a_14632_4688# VSS sg13_lv_nmos ad=0.14875p pd=1.16u as=0.187p ps=1.78u w=0.55u l=0.13u
x1246 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1247 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1248 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1249 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1250 a_15409_13743# a_14949_13701# a_15051_13844# VSS sg13_lv_nmos ad=0.31732p pd=1.805u as=0.2516p ps=2.16u w=0.74u l=0.13u
x1251 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1252 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1253 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1254 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1255 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1256 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1257 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1258 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1259 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1260 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1261 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1262 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1263 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1264 a_14758_15247# sg13_inv_1_0.Y VSS VSS sg13_lv_nmos ad=37.8f pd=0.6u as=0.1701p ps=1.65u w=0.42u l=0.13u
x1265 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1266 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1267 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1268 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1269 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1270 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1271 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1272 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1273 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1274 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1275 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1276 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1277 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1278 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1279 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1280 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1281 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1282 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1283 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1284 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1285 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1286 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1287 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1288 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1289 a_15801_16119# a_14859_16007# a_15599_16357# VDD sg13_lv_pmos ad=93.45f pd=0.865u as=0.2048p ps=1.63u w=0.42u l=0.13u
x1290 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1291 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1292 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1293 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1294 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1295 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1296 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1297 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1298 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1299 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1300 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1301 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1302 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1303 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1304 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1305 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1306 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1307 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1308 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1309 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1310 a_11076_16000# a_11050_15964# VSS VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.1626p ps=1.415u w=0.74u l=0.13u
x1311 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1312 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1313 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1314 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1315 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1316 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1317 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1318 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1319 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1320 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1321 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1322 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1323 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1324 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1325 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1326 a_11940_14040# a_12459_13844# a_13199_13799# VSS sg13_lv_nmos ad=0.3473p pd=2.71u as=0.12665p ps=1.145u w=0.74u l=0.13u
x1327 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1328 VDD sg13_inv_1_0.Y a_14506_15457# VDD sg13_lv_pmos ad=0.1563p pd=1.22u as=0.147p ps=1.54u w=0.42u l=0.13u
x1329 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1330 a_14532_14040# a_14506_13945# VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0.36237p ps=2.605u w=1u l=0.13u
x1331 a_13499_15996# sg13_nor2_1_0.Y sg13_dfrbpq_1_4.D VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.3808p ps=2.92u w=1.12u l=0.13u
x1332 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1333 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1334 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1335 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1336 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1337 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1338 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1339 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1340 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1341 a_12228_14922# sg13_nor2b_1_0.Y a_12134_14922# VSS sg13_lv_nmos ad=60.89999f pd=0.71u as=0.1428p ps=1.52u w=0.42u l=0.13u
x1342 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1343 a_12612_17064# a_12586_16969# VSS VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.1626p ps=1.415u w=0.74u l=0.13u
x1344 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1345 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1346 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1347 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1348 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1349 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1350 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1351 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1352 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1353 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1354 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1355 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1356 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1357 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1358 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1359 tx_start a_14248_23556# VDD VDD sg13_lv_pmos ad=0.42p pd=2.99u as=0.2114p ps=1.54u w=1.12u l=0.13u
x1360 a_15791_13799# a_14949_13701# a_15697_13799# VSS sg13_lv_nmos ad=0.12665p pd=1.145u as=0.1428p ps=1.52u w=0.42u l=0.13u
x1361 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1362 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1363 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1364 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1365 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1366 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1367 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1368 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1369 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1370 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1371 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1372 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1373 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1374 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1375 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1376 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1377 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1378 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1379 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1380 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1381 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1382 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1383 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1384 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1385 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1386 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1387 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1388 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1389 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1390 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1391 VDD a_13679_14845# a_13936_14726# VDD sg13_lv_pmos ad=0.4659p pd=3.65u as=79.8f ps=0.8u w=0.42u l=0.13u
x1392 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1393 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1394 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1395 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1396 a_14628_16421# a_14859_16007# a_14314_15964# VSS sg13_lv_nmos ad=0.2373p pd=1.97u as=79.8f ps=0.8u w=0.42u l=0.13u
x1397 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1398 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1399 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1400 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1401 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1402 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1403 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1404 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1405 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1406 a_15217_15998# a_14757_16007# a_14859_16007# VDD sg13_lv_pmos ad=0.41165p pd=2.12u as=0.3864p ps=2.93u w=1.12u l=0.13u
x1407 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1408 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1409 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1410 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1411 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1412 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1413 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1414 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1415 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1416 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1417 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1418 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1419 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1420 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1421 a_11914_13945# a_12357_13701# a_11654_13722# VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0.1296p ps=1.52u w=0.42u l=0.13u
x1422 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1423 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1424 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1425 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1426 a_11940_14040# a_11914_13945# VSS VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.1626p ps=1.415u w=0.74u l=0.13u
x1427 a_14820_13735# a_15051_13844# a_14506_13945# VSS sg13_lv_nmos ad=0.2373p pd=1.97u as=79.8f ps=0.8u w=0.42u l=0.13u
x1428 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1429 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1430 a_14949_13701# sg13_dfrbpq_1_0.CLK a_15409_14018# VDD sg13_lv_pmos ad=0.4088p pd=2.97u as=0.41165p ps=2.12u w=1.12u l=0.13u
x1431 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1432 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1433 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1434 VDD a_13199_13799# a_13456_13942# VDD sg13_lv_pmos ad=0.4659p pd=3.65u as=79.8f ps=0.8u w=0.42u l=0.13u
x1435 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1436 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1437 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1438 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1439 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1440 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1441 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1442 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1443 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1444 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1445 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1446 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1447 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1448 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1449 VDD sg13_buf_1_0.A a_13576_4688# VDD sg13_lv_pmos ad=0.2114p pd=1.54u as=0.2856p ps=2.36u w=0.84u l=0.13u
x1450 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1451 a_14128_16966# sg13_inv_1_0.Y a_14188_17061# VDD sg13_lv_pmos ad=79.8f pd=0.8u as=0.204p ps=1.835u w=0.42u l=0.13u
x1452 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1453 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1454 VDD clk a_7816_15996# VDD sg13_lv_pmos ad=0.2114p pd=1.54u as=0.2856p ps=2.36u w=0.84u l=0.13u
x1455 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1456 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1457 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1458 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1459 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1460 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1461 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1462 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1463 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1464 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1465 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1466 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1467 sg13_o21ai_1_0.A1 sg13_dfrbpq_1_5.Q VSS VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.2516p ps=2.16u w=0.74u l=0.13u
x1468 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1469 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1470 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1471 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1472 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1473 VSS sg13_inv_2_1.A a_17006_16388# VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=96.2f ps=1u w=0.74u l=0.13u
x1474 a_12817_13743# a_12357_13701# a_12459_13844# VSS sg13_lv_nmos ad=0.31732p pd=1.805u as=0.2516p ps=2.16u w=0.74u l=0.13u
x1475 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1476 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1477 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1478 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1479 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1480 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1481 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1482 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1483 sg13_buf_1_4.A a_13866_14020# VDD VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
x1484 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1485 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1486 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1487 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1488 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1489 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1490 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1491 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1492 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1493 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1494 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1495 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1496 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1497 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1498 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1499 VDD a_13679_14845# a_14346_14484# VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.3864p ps=2.93u w=1.12u l=0.13u
x1500 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1501 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1502 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1503 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1504 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1505 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1506 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1507 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1508 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1509 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1510 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1511 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1512 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1513 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1514 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1515 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1516 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1517 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1518 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1519 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1520 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1521 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1522 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1523 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1524 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1525 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1526 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1527 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1528 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1529 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1530 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1531 a_14532_14040# a_15051_13844# a_15791_13799# VSS sg13_lv_nmos ad=0.3473p pd=2.71u as=0.12665p ps=1.145u w=0.74u l=0.13u
x1532 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1533 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1534 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1535 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1536 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1537 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1538 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1539 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1540 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1541 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1542 VDD sg13_buf_1_0.A a_14248_4688# VDD sg13_lv_pmos ad=0.2114p pd=1.54u as=0.2856p ps=2.36u w=0.84u l=0.13u
x1543 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1544 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1545 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1546 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1547 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1548 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1549 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1550 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1551 a_13489_16767# a_13029_16725# a_13131_16868# VSS sg13_lv_nmos ad=0.31732p pd=1.805u as=0.2516p ps=2.16u w=0.74u l=0.13u
x1552 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1553 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1554 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1555 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1556 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1557 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1558 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1559 a_11940_14040# a_11914_13945# VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0.36237p ps=2.605u w=1u l=0.13u
x1560 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1561 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1562 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1563 VDD sg13_inv_1_0.Y a_14314_15964# VDD sg13_lv_pmos ad=0.1563p pd=1.22u as=0.147p ps=1.54u w=0.42u l=0.13u
x1564 VSS a_13679_14845# a_14346_14484# VSS sg13_lv_nmos ad=0.1406p pd=1.12u as=0.2516p ps=2.16u w=0.74u l=0.13u
x1565 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1566 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1567 VDD timer_done a_14152_10736# VDD sg13_lv_pmos ad=0.2114p pd=1.54u as=0.2856p ps=2.36u w=0.84u l=0.13u
x1568 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1569 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1570 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1571 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1572 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1573 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1574 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1575 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1576 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1577 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1578 sg13_dfrbpq_1_0.CLK a_7816_15996# VSS VSS sg13_lv_nmos ad=0.2886p pd=2.26u as=0.14875p ps=1.16u w=0.74u l=0.13u
x1579 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1580 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1581 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1582 a_12652_16119# a_12592_16238# a_12537_16119# VDD sg13_lv_pmos ad=0.204p pd=1.835u as=93.45f ps=0.865u w=0.42u l=0.13u
x1583 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1584 VSS sg13_a21o_1_0.A2 a_13838_12256# VSS sg13_lv_nmos ad=0.2176p pd=1.96u as=81.6f ps=0.895u w=0.64u l=0.13u
x1585 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1586 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1587 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1588 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1589 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1590 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1591 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1592 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1593 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1594 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1595 a_16294_14484# sg13_dfrbpq_1_1.Q a_16051_14746# VDD sg13_lv_pmos ad=0.2125p pd=1.425u as=0.35p ps=2.7u w=1u l=0.13u
x1596 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1597 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1598 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1599 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1600 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1601 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1602 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1603 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1604 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1605 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1606 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1607 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1608 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1609 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1610 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1611 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1612 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1613 sg13_dfrbpq_1_5.Q a_16266_15996# VSS VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.1406p ps=1.12u w=0.74u l=0.13u
x1614 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1615 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1616 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1617 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1618 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1619 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1620 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1621 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1622 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1623 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1624 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1625 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1626 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1627 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1628 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1629 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1630 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1631 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1632 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1633 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1634 a_14506_13945# a_14949_13701# a_14246_13722# VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0.1296p ps=1.52u w=0.42u l=0.13u
x1635 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1636 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1637 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1638 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1639 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1640 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1641 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1642 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1643 a_14820_13735# a_14532_14040# a_14758_13735# VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=37.8f ps=0.6u w=0.42u l=0.13u
x1644 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1645 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1646 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1647 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1648 a_12166_13735# sg13_inv_1_0.Y VSS VSS sg13_lv_nmos ad=37.8f pd=0.6u as=0.1701p ps=1.65u w=0.42u l=0.13u
x1649 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1650 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1651 a_12357_13701# sg13_dfrbpq_1_0.CLK a_12817_14018# VDD sg13_lv_pmos ad=0.4088p pd=2.97u as=0.41165p ps=2.12u w=1.12u l=0.13u
x1652 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1653 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1654 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1655 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1656 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1657 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1658 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1659 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1660 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1661 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1662 VSS sg13_a21o_1_1.A2 a_16430_14832# VSS sg13_lv_nmos ad=0.2176p pd=1.96u as=81.6f ps=0.895u w=0.64u l=0.13u
x1663 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1664 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1665 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1666 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1667 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1668 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1669 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1670 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1671 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1672 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1673 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1674 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1675 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1676 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1677 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1678 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1679 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1680 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1681 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1682 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1683 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1684 VSS sg13_buf_1_0.A a_13576_4688# VSS sg13_lv_nmos ad=0.14875p pd=1.16u as=0.187p ps=1.78u w=0.55u l=0.13u
x1685 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1686 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1687 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1688 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1689 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1690 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1691 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1692 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1693 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1694 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1695 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1696 sg13_dfrbpq_1_1.Q a_16458_14020# VDD VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
x1697 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1698 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1699 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1700 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1701 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1702 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1703 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1704 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1705 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1706 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1707 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1708 sg13_inv_1_1.A sg13_dfrbpq_1_5.Q a_16735_15972# VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2716p ps=1.605u w=1.12u l=0.13u
x1709 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1710 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1711 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1712 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1713 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1714 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1715 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1716 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1717 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1718 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1719 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1720 a_14949_15213# sg13_dfrbpq_1_0.CLK a_15409_15255# VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.31732p ps=1.805u w=0.74u l=0.13u
x1721 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1722 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1723 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1724 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1725 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1726 VSS sg13_buf_1_5.X sg13_a21o_1_0.A2 VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.1406p ps=1.12u w=0.74u l=0.13u
x1727 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1728 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1729 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1730 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1731 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1732 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1733 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1734 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1735 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1736 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1737 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1738 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1739 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1740 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1741 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1742 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1743 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1744 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1745 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1746 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1747 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1748 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1749 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1750 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1751 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1752 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1753 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1754 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1755 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1756 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1757 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1758 a_12754_16434# sg13_inv_1_0.Y VSS VSS sg13_lv_nmos ad=37.8f pd=0.6u as=79.8f ps=0.8u w=0.42u l=0.13u
x1759 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1760 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1761 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1762 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1763 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1764 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1765 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1766 VDD sg13_buf_1_4.A a_13702_12532# VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0.2125p ps=1.425u w=1u l=0.13u
x1767 a_11493_16007# sg13_dfrbpq_1_0.CLK a_11953_15998# VDD sg13_lv_pmos ad=0.4088p pd=2.97u as=0.41165p ps=2.12u w=1.12u l=0.13u
x1768 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1769 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1770 a_16210_13722# sg13_inv_1_0.Y VSS VSS sg13_lv_nmos ad=37.8f pd=0.6u as=79.8f ps=0.8u w=0.42u l=0.13u
x1771 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1772 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1773 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1774 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1775 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1776 VSS sg13_buf_1_0.A a_14248_4688# VSS sg13_lv_nmos ad=0.14875p pd=1.16u as=0.187p ps=1.78u w=0.55u l=0.13u
x1777 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1778 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1779 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1780 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1781 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1782 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1783 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1784 sg13_buf_1_5.X a_14152_10736# VDD VDD sg13_lv_pmos ad=0.42p pd=2.99u as=0.2114p ps=1.54u w=1.12u l=0.13u
x1785 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1786 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1787 a_14949_15213# sg13_dfrbpq_1_0.CLK a_15409_15530# VDD sg13_lv_pmos ad=0.4088p pd=2.97u as=0.41165p ps=2.12u w=1.12u l=0.13u
x1788 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1789 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1790 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1791 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1792 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1793 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1794 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1795 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1796 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1797 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1798 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1799 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1800 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1801 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1802 sg13_and2_1_0.X a_14061_12256# VSS VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.1331p ps=1.12u w=0.74u l=0.13u
x1803 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1804 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1805 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1806 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1807 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1808 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1809 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1810 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1811 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1812 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1813 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1814 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1815 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1816 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1817 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1818 a_13489_17042# a_13029_16725# a_13131_16868# VDD sg13_lv_pmos ad=0.41165p pd=2.12u as=0.3864p ps=2.93u w=1.12u l=0.13u
x1819 a_15856_16238# a_15599_16357# a_16018_16434# VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=37.8f ps=0.6u w=0.42u l=0.13u
x1820 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1821 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1822 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1823 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1824 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1825 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1826 a_10790_16434# a_11595_16007# a_11050_15964# VDD sg13_lv_pmos ad=0.1428p pd=1.52u as=79.8f ps=0.8u w=0.42u l=0.13u
x1827 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1828 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1829 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1830 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1831 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1832 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1833 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1834 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1835 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1836 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1837 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1838 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1839 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1840 a_12612_17064# a_13131_16868# a_13871_16823# VSS sg13_lv_nmos ad=0.3473p pd=2.71u as=0.12665p ps=1.145u w=0.74u l=0.13u
x1841 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1842 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1843 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1844 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1845 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1846 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1847 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1848 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1849 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1850 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1851 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1852 Timer_en a_13768_10736# VSS VSS sg13_lv_nmos ad=0.2886p pd=2.26u as=0.14875p ps=1.16u w=0.74u l=0.13u
x1853 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1854 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1855 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1856 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1857 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1858 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1859 a_16430_14832# sg13_dfrbpq_1_3.Q a_16051_14746# VSS sg13_lv_nmos ad=81.6f pd=0.895u as=0.1216p ps=1.02u w=0.64u l=0.13u
x1860 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1861 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1862 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1863 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1864 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1865 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1866 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1867 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1868 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1869 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1870 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1871 VDD sg13_buf_1_0.A a_14440_5412# VDD sg13_lv_pmos ad=0.2114p pd=1.54u as=0.2856p ps=2.36u w=0.84u l=0.13u
x1872 a_14155_12256# sg13_buf_1_4.A a_14061_12256# VSS sg13_lv_nmos ad=0.1216p pd=1.02u as=0.2176p ps=1.96u w=0.64u l=0.13u
x1873 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1874 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1875 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1876 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1877 a_14246_15234# a_15051_15356# a_14506_15457# VDD sg13_lv_pmos ad=0.1428p pd=1.52u as=79.8f ps=0.8u w=0.42u l=0.13u
x1878 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1879 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1880 a_14758_13735# sg13_inv_1_0.Y VSS VSS sg13_lv_nmos ad=37.8f pd=0.6u as=0.1701p ps=1.65u w=0.42u l=0.13u
x1881 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1882 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1883 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1884 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1885 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1886 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1887 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1888 a_16108_15549# a_16048_15454# a_15993_15549# VDD sg13_lv_pmos ad=0.204p pd=1.835u as=93.45f ps=0.865u w=0.42u l=0.13u
x1889 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1890 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1891 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1892 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1893 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1894 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1895 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1896 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1897 a_13871_16823# a_13029_16725# a_13777_16823# VSS sg13_lv_nmos ad=0.12665p pd=1.145u as=0.1428p ps=1.52u w=0.42u l=0.13u
x1898 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1899 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1900 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1901 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1902 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1903 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1904 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1905 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1906 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1907 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1908 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1909 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1910 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1911 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1912 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1913 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1914 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1915 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1916 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1917 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1918 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1919 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1920 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1921 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1922 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1923 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1924 VDD sg13_inv_1_0.Y a_11914_13945# VDD sg13_lv_pmos ad=0.1563p pd=1.22u as=0.147p ps=1.54u w=0.42u l=0.13u
x1925 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1926 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1927 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1928 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1929 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1930 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1931 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1932 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1933 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1934 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1935 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1936 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1937 VSS a_15791_15311# a_16458_15532# VSS sg13_lv_nmos ad=0.1406p pd=1.12u as=0.2516p ps=2.16u w=0.74u l=0.13u
x1938 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1939 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1940 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1941 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1942 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1943 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1944 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1945 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1946 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1947 a_12134_14922# a_12939_14495# a_12394_14452# VDD sg13_lv_pmos ad=0.1428p pd=1.52u as=79.8f ps=0.8u w=0.42u l=0.13u
x1948 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1949 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1950 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1951 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1952 a_12900_16759# a_12612_17064# a_12838_16759# VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=37.8f ps=0.6u w=0.42u l=0.13u
x1953 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1954 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1955 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1956 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1957 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1958 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1959 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1960 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1961 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1962 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1963 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1964 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1965 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1966 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1967 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1968 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1969 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1970 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1971 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1972 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1973 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1974 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1975 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1976 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1977 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1978 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1979 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1980 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1981 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1982 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1983 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1984 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1985 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1986 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1987 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1988 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1989 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1990 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1991 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x1992 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1993 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x1994 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1995 sg13_a21oi_1_0.A1 a_14538_17044# VDD VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
x1996 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x1997 VDD sg13_nor2_1_0.A a_12046_15276# VDD sg13_lv_pmos ad=0.2618p pd=1.63u as=0.2856p ps=2.36u w=0.84u l=0.13u
x1998 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x1999 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2000 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2001 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2002 a_13618_13722# sg13_inv_1_0.Y VSS VSS sg13_lv_nmos ad=37.8f pd=0.6u as=79.8f ps=0.8u w=0.42u l=0.13u
x2003 VDD sg13_a21oi_1_0.A2 a_14235_17564# VDD sg13_lv_pmos ad=0.2198p pd=1.53u as=0.2856p ps=2.36u w=0.84u l=0.13u
x2004 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2005 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2006 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2007 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2008 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2009 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2010 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2011 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2012 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2013 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2014 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2015 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2016 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2017 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2018 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2019 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2020 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2021 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2022 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2023 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2024 a_14340_16000# a_14314_15964# VSS VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.1626p ps=1.415u w=0.74u l=0.13u
x2025 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2026 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2027 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2028 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2029 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2030 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2031 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2032 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2033 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2034 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2035 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2036 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2037 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2038 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2039 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2040 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2041 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2042 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2043 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2044 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2045 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2046 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2047 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2048 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2049 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2050 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2051 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2052 sg13_nor2b_1_0.Y sg13_nor2_1_0.B a_12268_15532# VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.1176p ps=1.33u w=1.12u l=0.13u
x2053 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2054 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2055 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2056 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2057 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2058 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2059 sg13_a21o_1_1.A2 sg13_inv_2_1.A VSS VSS sg13_lv_nmos ad=0.1406p pd=1.12u as=0.2516p ps=2.16u w=0.74u l=0.13u
x2060 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2061 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2062 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2063 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2064 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2065 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2066 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2067 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2068 a_14506_15457# a_14949_15213# a_14889_15625# VDD sg13_lv_pmos ad=79.8f pd=0.8u as=63f ps=0.72u w=0.42u l=0.13u
x2069 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2070 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2071 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2072 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2073 a_14290_16746# sg13_inv_1_0.Y VSS VSS sg13_lv_nmos ad=37.8f pd=0.6u as=79.8f ps=0.8u w=0.42u l=0.13u
x2074 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2075 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2076 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2077 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2078 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2079 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2080 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2081 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2082 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2083 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2084 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2085 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2086 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2087 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2088 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2089 VSS sg13_nor2_1_0.B sg13_nor2b_1_0.Y VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.1406p ps=1.12u w=0.74u l=0.13u
x2090 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2091 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2092 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2093 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2094 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2095 VSS sg13_buf_1_5.X a_14155_12256# VSS sg13_lv_nmos ad=0.1331p pd=1.12u as=0.1216p ps=1.02u w=0.64u l=0.13u
x2096 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2097 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2098 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2099 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2100 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2101 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2102 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2103 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2104 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2105 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2106 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2107 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2108 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2109 VSS sg13_nor2_1_0.A a_12046_15276# VSS sg13_lv_nmos ad=0.17255p pd=1.25u as=0.187p ps=1.78u w=0.55u l=0.13u
x2110 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2111 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2112 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2113 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2114 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2115 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2116 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2117 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2118 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2119 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2120 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2121 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2122 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2123 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2124 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2125 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2126 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2127 VDD sg13_inv_1_0.Y a_14506_13945# VDD sg13_lv_pmos ad=0.1563p pd=1.22u as=0.147p ps=1.54u w=0.42u l=0.13u
x2128 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2129 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2130 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2131 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2132 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2133 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2134 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2135 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2136 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2137 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2138 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2139 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2140 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2141 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2142 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2143 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2144 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2145 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2146 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2147 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2148 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2149 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2150 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2151 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2152 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2153 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2154 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2155 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2156 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2157 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2158 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2159 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2160 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2161 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2162 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2163 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2164 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2165 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2166 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2167 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2168 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2169 a_12838_16759# sg13_inv_1_0.Y VSS VSS sg13_lv_nmos ad=37.8f pd=0.6u as=0.1701p ps=1.65u w=0.42u l=0.13u
x2170 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2171 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2172 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2173 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2174 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2175 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2176 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2177 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2178 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2179 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2180 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2181 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2182 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2183 a_15599_16357# a_14757_16007# a_15505_16357# VSS sg13_lv_nmos ad=0.12665p pd=1.145u as=0.1428p ps=1.52u w=0.42u l=0.13u
x2184 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2185 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2186 a_15856_16238# sg13_inv_1_0.Y a_15916_16119# VDD sg13_lv_pmos ad=79.8f pd=0.8u as=0.204p ps=1.835u w=0.42u l=0.13u
x2187 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2188 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2189 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2190 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2191 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2192 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2193 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2194 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2195 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2196 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2197 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2198 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2199 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2200 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2201 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2202 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2203 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2204 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2205 VDD sg13_dfrbpq_1_1.Q a_17128_13760# VDD sg13_lv_pmos ad=0.2114p pd=1.54u as=0.2856p ps=2.36u w=0.84u l=0.13u
x2206 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2207 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2208 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2209 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2210 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2211 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2212 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2213 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2214 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2215 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2216 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2217 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2218 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2219 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2220 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2221 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2222 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2223 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2224 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2225 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2226 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2227 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2228 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2229 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2230 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2231 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2232 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2233 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2234 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2235 a_15791_15311# a_14949_15213# a_14532_15552# VDD sg13_lv_pmos ad=0.2048p pd=1.63u as=0.34p ps=2.68u w=1u l=0.13u
x2236 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2237 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2238 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2239 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2240 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2241 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2242 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2243 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2244 a_16048_15454# a_15791_15311# a_16210_15234# VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=37.8f ps=0.6u w=0.42u l=0.13u
x2245 VSS a_13936_14726# a_13585_14845# VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
x2246 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2247 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2248 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2249 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2250 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2251 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2252 VDD wake_up_sg a_10024_15996# VDD sg13_lv_pmos ad=0.2114p pd=1.54u as=0.2856p ps=2.36u w=0.84u l=0.13u
x2253 sg13_a21o_1_0.A2 sg13_buf_1_5.X VDD VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.3808p ps=2.92u w=1.12u l=0.13u
x2254 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2255 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2256 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2257 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2258 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2259 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2260 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2261 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2262 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2263 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2264 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2265 a_12777_14531# a_12420_14488# VDD VDD sg13_lv_pmos ad=63f pd=0.72u as=0.1563p ps=1.22u w=0.42u l=0.13u
x2266 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2267 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2268 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2269 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2270 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2271 a_12134_14922# sg13_nor2b_1_0.Y VDD VDD sg13_lv_pmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
x2272 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2273 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2274 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2275 sg13_nor2_1_0.A a_10024_15996# VDD VDD sg13_lv_pmos ad=0.42p pd=2.99u as=0.2114p ps=1.54u w=1.12u l=0.13u
x2276 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2277 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2278 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2279 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2280 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2281 a_14314_15964# a_14757_16007# a_14697_16043# VDD sg13_lv_pmos ad=79.8f pd=0.8u as=63f ps=0.72u w=0.42u l=0.13u
x2282 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2283 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2284 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2285 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2286 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2287 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2288 sg13_a21o_1_1.A2 sg13_inv_2_1.A VDD VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.3808p ps=2.92u w=1.12u l=0.13u
x2289 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2290 a_14061_12256# sg13_buf_1_4.A VDD VDD sg13_lv_pmos ad=0.1596p pd=1.22u as=0.2856p ps=2.36u w=0.84u l=0.13u
x2291 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2292 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2293 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2294 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2295 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2296 sg13_inv_2_1.A a_17800_15272# VSS VSS sg13_lv_nmos ad=0.2886p pd=2.26u as=0.14875p ps=1.16u w=0.74u l=0.13u
x2297 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2298 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2299 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2300 adc_start a_17128_13760# VSS VSS sg13_lv_nmos ad=0.2886p pd=2.26u as=0.14875p ps=1.16u w=0.74u l=0.13u
x2301 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2302 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2303 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2304 a_14949_13701# sg13_dfrbpq_1_0.CLK a_15409_13743# VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.31732p ps=1.805u w=0.74u l=0.13u
x2305 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2306 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2307 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2308 a_14998_16742# sg13_a22oi_1_0.B2 VSS VSS sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.15u
x2309 a_11076_16000# a_11050_15964# VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0.36237p ps=2.605u w=1u l=0.13u
x2310 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2311 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2312 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2313 a_11302_16421# sg13_inv_1_0.Y VSS VSS sg13_lv_nmos ad=37.8f pd=0.6u as=0.1701p ps=1.65u w=0.42u l=0.13u
x2314 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2315 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2316 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2317 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2318 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2319 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2320 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2321 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2322 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2323 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2324 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2325 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2326 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2327 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2328 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2329 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2330 sg13_a22oi_1_0.B2 a_15976_25068# VSS VSS sg13_lv_nmos ad=0.2886p pd=2.26u as=0.14875p ps=1.16u w=0.74u l=0.13u
x2331 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2332 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2333 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2334 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2335 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2336 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2337 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2338 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2339 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2340 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2341 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2342 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2343 VSS sg13_a21oi_1_0.A2 a_13601_16344# VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.1406p ps=1.12u w=0.74u l=0.13u
x2344 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2345 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2346 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2347 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2348 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2349 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2350 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2351 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2352 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2353 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2354 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2355 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2356 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2357 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2358 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2359 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2360 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2361 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2362 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2363 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2364 a_11050_15964# a_11493_16007# a_10790_16434# VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0.1296p ps=1.52u w=0.42u l=0.13u
x2365 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2366 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2367 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2368 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2369 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2370 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2371 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2372 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2373 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2374 VSS sg13_a21oi_1_0.A2 a_14235_17564# VSS sg13_lv_nmos ad=0.14505p pd=1.15u as=0.187p ps=1.78u w=0.55u l=0.13u
x2375 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2376 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2377 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2378 sg13_nor2_1_0.B a_13002_15996# VDD VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
x2379 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2380 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2381 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2382 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2383 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2384 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2385 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2386 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2387 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2388 a_12326_16746# sg13_dfrbpq_1_6.D VDD VDD sg13_lv_pmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
x2389 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2390 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2391 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2392 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2393 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2394 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2395 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2396 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2397 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2398 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2399 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2400 a_13297_14837# a_12837_14495# a_12939_14495# VSS sg13_lv_nmos ad=0.31732p pd=1.805u as=0.2516p ps=2.16u w=0.74u l=0.13u
x2401 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2402 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2403 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2404 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2405 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2406 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2407 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2408 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2409 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2410 VDD uart_busy a_15976_25068# VDD sg13_lv_pmos ad=0.2114p pd=1.54u as=0.2856p ps=2.36u w=0.84u l=0.13u
x2411 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2412 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2413 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2414 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2415 sg13_a21oi_1_0.A2 a_13960_25068# VDD VDD sg13_lv_pmos ad=0.42p pd=2.99u as=0.2114p ps=1.54u w=1.12u l=0.13u
x2416 VSS sg13_inv_1_0.Y a_10884_16434# VSS sg13_lv_nmos ad=0.1626p pd=1.415u as=60.89999f ps=0.71u w=0.42u l=0.13u
x2417 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2418 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2419 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2420 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2421 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2422 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2423 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2424 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2425 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2426 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2427 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2428 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2429 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2430 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2431 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2432 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2433 a_11953_15998# a_11493_16007# a_11595_16007# VDD sg13_lv_pmos ad=0.41165p pd=2.12u as=0.3864p ps=2.93u w=1.12u l=0.13u
x2434 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2435 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2436 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2437 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2438 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2439 a_12335_16357# a_11493_16007# a_11076_16000# VDD sg13_lv_pmos ad=0.2048p pd=1.63u as=0.34p ps=2.68u w=1u l=0.13u
x2440 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2441 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2442 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2443 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2444 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2445 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2446 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2447 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2448 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2449 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2450 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2451 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2452 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2453 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2454 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2455 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2456 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2457 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2458 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2459 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2460 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2461 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2462 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2463 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2464 a_14757_16007# sg13_dfrbpq_1_0.CLK a_15217_15998# VDD sg13_lv_pmos ad=0.4088p pd=2.97u as=0.41165p ps=2.12u w=1.12u l=0.13u
x2465 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2466 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2467 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2468 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2469 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2470 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2471 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2472 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2473 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2474 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2475 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2476 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2477 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2478 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2479 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2480 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2481 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2482 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2483 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2484 a_12394_14452# a_12837_14495# a_12134_14922# VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0.1296p ps=1.52u w=0.42u l=0.13u
x2485 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2486 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2487 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2488 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2489 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2490 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2491 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2492 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2493 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2494 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2495 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2496 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2497 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2498 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2499 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2500 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2501 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2502 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2503 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2504 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2505 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2506 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2507 VSS a_13459_12404# sg13_a21o_1_0.X VSS sg13_lv_nmos ad=0.15745p pd=1.175u as=0.2351p ps=2.16u w=0.74u l=0.13u
x2508 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2509 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2510 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2511 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2512 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2513 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2514 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2515 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2516 a_13679_14845# a_12837_14495# a_12420_14488# VDD sg13_lv_pmos ad=0.2048p pd=1.63u as=0.34p ps=2.68u w=1u l=0.13u
x2517 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2518 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2519 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2520 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2521 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2522 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2523 VSS a_15791_13799# a_16458_14020# VSS sg13_lv_nmos ad=0.1406p pd=1.12u as=0.2516p ps=2.16u w=0.74u l=0.13u
x2524 VDD sg13_a21oi_1_0.A1 a_13499_15996# VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
x2525 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2526 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2527 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2528 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2529 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2530 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2531 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2532 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2533 VDD sg13_buf_1_5.X a_14061_12256# VDD sg13_lv_pmos ad=0.1918p pd=1.5u as=0.1596p ps=1.22u w=0.84u l=0.13u
x2534 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2535 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2536 a_12357_13701# sg13_dfrbpq_1_0.CLK a_12817_13743# VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.31732p ps=1.805u w=0.74u l=0.13u
x2537 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2538 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2539 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2540 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2541 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2542 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2543 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2544 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2545 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2546 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2547 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2548 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2549 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2550 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2551 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2552 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2553 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2554 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2555 VSS sg13_buf_1_4.A a_13768_10736# VSS sg13_lv_nmos ad=0.14875p pd=1.16u as=0.187p ps=1.78u w=0.55u l=0.13u
x2556 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2557 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2558 tx_start a_14248_23556# VSS VSS sg13_lv_nmos ad=0.2886p pd=2.26u as=0.14875p ps=1.16u w=0.74u l=0.13u
x2559 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2560 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2561 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2562 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2563 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2564 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2565 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2566 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2567 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2568 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2569 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2570 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2571 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2572 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2573 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2574 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2575 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2576 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2577 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2578 VSS a_12335_16357# a_13002_15996# VSS sg13_lv_nmos ad=0.1406p pd=1.12u as=0.2516p ps=2.16u w=0.74u l=0.13u
x2579 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2580 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2581 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2582 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2583 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2584 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2585 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2586 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2587 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2588 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2589 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2590 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2591 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2592 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2593 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2594 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2595 a_14246_15234# sg13_dfrbpq_1_3.D VDD VDD sg13_lv_pmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
x2596 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2597 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2598 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2599 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2600 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2601 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2602 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2603 a_13029_16725# sg13_dfrbpq_1_0.CLK a_13489_16767# VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.31732p ps=1.805u w=0.74u l=0.13u
x2604 a_15993_15549# a_15051_15356# a_15791_15311# VDD sg13_lv_pmos ad=93.45f pd=0.865u as=0.2048p ps=1.63u w=0.42u l=0.13u
x2605 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2606 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2607 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2608 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2609 a_10884_16434# sg13_dfrbpq_1_4.D a_10790_16434# VSS sg13_lv_nmos ad=60.89999f pd=0.71u as=0.1428p ps=1.52u w=0.42u l=0.13u
x2610 a_12228_13735# a_12459_13844# a_11914_13945# VSS sg13_lv_nmos ad=0.2373p pd=1.97u as=79.8f ps=0.8u w=0.42u l=0.13u
x2611 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2612 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2613 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2614 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2615 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2616 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2617 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2618 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2619 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2620 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2621 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2622 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2623 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2624 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2625 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2626 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2627 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2628 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2629 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2630 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2631 a_16735_16388# sg13_dfrbpq_1_5.Q VSS VSS sg13_lv_nmos ad=0.13875p pd=1.115u as=0.2553p ps=2.17u w=0.74u l=0.13u
x2632 VDD sg13_a21oi_1_0.A1 a_14248_23556# VDD sg13_lv_pmos ad=0.2114p pd=1.54u as=0.2856p ps=2.36u w=0.84u l=0.13u
x2633 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2634 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2635 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2636 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2637 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2638 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2639 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2640 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2641 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2642 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2643 VDD a_13871_16823# a_14128_16966# VDD sg13_lv_pmos ad=0.4659p pd=3.65u as=79.8f ps=0.8u w=0.42u l=0.13u
x2644 a_11914_13945# a_12357_13701# a_12297_14113# VDD sg13_lv_pmos ad=79.8f pd=0.8u as=63f ps=0.72u w=0.42u l=0.13u
x2645 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2646 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2647 VSS sg13_dfrbpq_1_1.Q a_17128_13760# VSS sg13_lv_nmos ad=0.14875p pd=1.16u as=0.187p ps=1.78u w=0.55u l=0.13u
x2648 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2649 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2650 a_14246_13722# a_15051_13844# a_14506_13945# VDD sg13_lv_pmos ad=0.1428p pd=1.52u as=79.8f ps=0.8u w=0.42u l=0.13u
x2651 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2652 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2653 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2654 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2655 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2656 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2657 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2658 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2659 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2660 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2661 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2662 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2663 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2664 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2665 a_16108_14037# a_16048_13942# a_15993_14037# VDD sg13_lv_pmos ad=0.204p pd=1.835u as=93.45f ps=0.865u w=0.42u l=0.13u
x2666 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2667 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2668 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2669 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2670 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2671 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2672 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2673 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2674 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2675 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2676 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2677 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2678 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2679 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2680 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2681 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2682 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2683 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2684 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2685 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2686 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2687 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2688 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2689 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2690 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2691 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2692 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2693 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2694 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2695 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2696 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2697 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2698 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2699 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2700 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2701 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2702 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2703 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2704 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2705 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2706 sg13_buf_1_0.A a_14346_14484# VDD VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
x2707 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2708 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2709 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2710 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2711 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2712 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2713 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2714 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2715 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2716 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2717 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2718 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2719 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2720 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2721 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2722 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2723 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2724 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2725 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2726 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2727 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2728 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2729 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2730 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2731 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2732 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2733 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2734 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2735 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2736 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2737 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2738 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2739 a_12586_16969# a_13029_16725# a_12969_17137# VDD sg13_lv_pmos ad=79.8f pd=0.8u as=63f ps=0.72u w=0.42u l=0.13u
x2740 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2741 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2742 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2743 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2744 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2745 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2746 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2747 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2748 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2749 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2750 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2751 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2752 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2753 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2754 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2755 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2756 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2757 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2758 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2759 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2760 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2761 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2762 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2763 a_12228_13735# a_11940_14040# a_12166_13735# VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=37.8f ps=0.6u w=0.42u l=0.13u
x2764 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2765 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2766 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2767 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2768 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2769 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2770 VSS a_13199_13799# a_13866_14020# VSS sg13_lv_nmos ad=0.1406p pd=1.12u as=0.2516p ps=2.16u w=0.74u l=0.13u
x2771 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2772 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2773 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2774 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2775 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2776 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2777 sg13_nor2_1_0.Y sg13_nor2_1_0.B a_12650_15532# VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.1176p ps=1.33u w=1.12u l=0.13u
x2778 sg13_buf_1_0.A a_14346_14484# VSS VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.1406p ps=1.12u w=0.74u l=0.13u
x2779 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2780 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2781 sg13_dfrbpq_1_6.D sg13_o21ai_1_0.B1 a_14998_16742# VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.1406p ps=1.12u w=0.74u l=0.15u
x2782 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2783 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2784 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2785 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2786 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2787 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2788 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2789 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2790 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2791 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2792 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2793 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2794 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2795 a_12335_16357# a_11493_16007# a_12241_16357# VSS sg13_lv_nmos ad=0.12665p pd=1.145u as=0.1428p ps=1.52u w=0.42u l=0.13u
x2796 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2797 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2798 a_12592_16238# sg13_inv_1_0.Y a_12652_16119# VDD sg13_lv_pmos ad=79.8f pd=0.8u as=0.204p ps=1.835u w=0.42u l=0.13u
x2799 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2800 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2801 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2802 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2803 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2804 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2805 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2806 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2807 sg13_inv_1_1.Y sg13_inv_1_1.A VSS VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.2516p ps=2.16u w=0.74u l=0.13u
x2808 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2809 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2810 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2811 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2812 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2813 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2814 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2815 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2816 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2817 a_12420_14488# a_12939_14495# a_13679_14845# VSS sg13_lv_nmos ad=0.3473p pd=2.71u as=0.12665p ps=1.145u w=0.74u l=0.13u
x2818 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2819 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2820 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2821 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2822 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2823 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2824 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2825 VSS sg13_inv_1_0.Y a_14340_15234# VSS sg13_lv_nmos ad=0.1626p pd=1.415u as=60.89999f ps=0.71u w=0.42u l=0.13u
x2826 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2827 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2828 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2829 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2830 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2831 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2832 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2833 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2834 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2835 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2836 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2837 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2838 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2839 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2840 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2841 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2842 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2843 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2844 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2845 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2846 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2847 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2848 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2849 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2850 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2851 VSS a_13871_16823# a_14538_17044# VSS sg13_lv_nmos ad=0.1406p pd=1.12u as=0.2516p ps=2.16u w=0.74u l=0.13u
x2852 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2853 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2854 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2855 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2856 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2857 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2858 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2859 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2860 a_13199_13799# a_12357_13701# a_11940_14040# VDD sg13_lv_pmos ad=0.2048p pd=1.63u as=0.34p ps=2.68u w=1u l=0.13u
x2861 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2862 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2863 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2864 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2865 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2866 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2867 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2868 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2869 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2870 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2871 VSS sg13_buf_1_0.A a_14440_5412# VSS sg13_lv_nmos ad=0.14875p pd=1.16u as=0.187p ps=1.78u w=0.55u l=0.13u
x2872 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2873 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2874 VSS sg13_o21ai_1_0.A1 a_14998_16742# VSS sg13_lv_nmos ad=0.1406p pd=1.12u as=0.2516p ps=2.16u w=0.74u l=0.15u
x2875 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2876 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2877 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2878 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2879 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2880 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2881 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2882 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2883 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2884 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2885 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2886 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2887 a_14506_13945# a_14949_13701# a_14889_14113# VDD sg13_lv_pmos ad=79.8f pd=0.8u as=63f ps=0.72u w=0.42u l=0.13u
x2888 a_16048_13942# a_15791_13799# a_16210_13722# VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=37.8f ps=0.6u w=0.42u l=0.13u
x2889 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2890 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2891 VSS clk a_7816_15996# VSS sg13_lv_nmos ad=0.14875p pd=1.16u as=0.187p ps=1.78u w=0.55u l=0.13u
x2892 VDD a_15599_16357# a_16266_15996# VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.3864p ps=2.93u w=1.12u l=0.13u
x2893 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2894 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2895 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2896 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2897 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2898 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2899 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2900 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2901 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2902 a_13029_16725# sg13_dfrbpq_1_0.CLK a_13489_17042# VDD sg13_lv_pmos ad=0.4088p pd=2.97u as=0.41165p ps=2.12u w=1.12u l=0.13u
x2903 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2904 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2905 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2906 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2907 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2908 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2909 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2910 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2911 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2912 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2913 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2914 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2915 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2916 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2917 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2918 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2919 a_13516_14037# a_13456_13942# a_13401_14037# VDD sg13_lv_pmos ad=0.204p pd=1.835u as=93.45f ps=0.865u w=0.42u l=0.13u
x2920 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2921 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2922 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2923 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2924 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2925 a_14148_16434# sg13_inv_1_1.Y a_14054_16434# VSS sg13_lv_nmos ad=60.89999f pd=0.71u as=0.1428p ps=1.52u w=0.42u l=0.13u
x2926 a_16735_15972# sg13_a22oi_1_0.B2 sg13_inv_1_1.A VDD sg13_lv_pmos ad=0.2744p pd=1.61u as=0.2128p ps=1.5u w=1.12u l=0.13u
x2927 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2928 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2929 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2930 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2931 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2932 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2933 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2934 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2935 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2936 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2937 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2938 sg13_nor2_1_0.Y sg13_nor2_1_0.A VSS VSS sg13_lv_nmos ad=0.1406p pd=1.12u as=0.2516p ps=2.16u w=0.74u l=0.13u
x2939 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2940 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2941 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2942 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2943 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2944 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2945 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2946 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2947 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2948 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2949 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2950 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2951 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2952 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2953 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2954 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2955 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2956 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2957 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2958 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2959 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2960 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2961 a_12420_16746# sg13_dfrbpq_1_6.D a_12326_16746# VSS sg13_lv_nmos ad=60.89999f pd=0.71u as=0.1428p ps=1.52u w=0.42u l=0.13u
x2962 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2963 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2964 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2965 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2966 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2967 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2968 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2969 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2970 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2971 VDD a_15599_16357# a_15856_16238# VDD sg13_lv_pmos ad=0.4659p pd=3.65u as=79.8f ps=0.8u w=0.42u l=0.13u
x2972 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2973 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2974 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2975 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2976 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2977 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2978 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2979 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2980 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2981 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2982 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2983 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2984 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2985 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2986 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x2987 a_12326_16746# a_13131_16868# a_12586_16969# VDD sg13_lv_pmos ad=0.1428p pd=1.52u as=79.8f ps=0.8u w=0.42u l=0.13u
x2988 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2989 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2990 a_13702_12532# sg13_a21o_1_0.A2 VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0.19p ps=1.38u w=1u l=0.13u
x2991 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2992 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2993 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2994 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2995 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2996 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x2997 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x2998 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x2999 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3000 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3001 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3002 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3003 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3004 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3005 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3006 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3007 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3008 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3009 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3010 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3011 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3012 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3013 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3014 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3015 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3016 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3017 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3018 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3019 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3020 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3021 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3022 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3023 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3024 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3025 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3026 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3027 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3028 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3029 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3030 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3031 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3032 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3033 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3034 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3035 VDD a_12335_16357# a_12592_16238# VDD sg13_lv_pmos ad=0.4659p pd=3.65u as=79.8f ps=0.8u w=0.42u l=0.13u
x3036 VDD sg13_dfrbpq_1_3.Q a_16294_14484# VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0.2125p ps=1.425u w=1u l=0.13u
x3037 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3038 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3039 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3040 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3041 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3042 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3043 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3044 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3045 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3046 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3047 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3048 a_14098_14922# sg13_inv_1_0.Y VSS VSS sg13_lv_nmos ad=37.8f pd=0.6u as=79.8f ps=0.8u w=0.42u l=0.13u
x3049 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3050 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3051 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3052 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3053 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3054 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3055 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3056 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3057 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3058 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3059 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3060 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3061 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3062 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3063 VDD sg13_buf_1_5.X sg13_a21o_1_0.A2 VDD sg13_lv_pmos ad=0.3864p pd=2.93u as=0.2128p ps=1.5u w=1.12u l=0.13u
x3064 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3065 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3066 a_14566_16421# sg13_inv_1_0.Y VSS VSS sg13_lv_nmos ad=37.8f pd=0.6u as=0.1701p ps=1.65u w=0.42u l=0.13u
x3067 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3068 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3069 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3070 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3071 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3072 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3073 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3074 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3075 a_15791_13799# a_14949_13701# a_14532_14040# VDD sg13_lv_pmos ad=0.2048p pd=1.63u as=0.34p ps=2.68u w=1u l=0.13u
x3076 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3077 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3078 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3079 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3080 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3081 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3082 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3083 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3084 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3085 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3086 sg13_buf_1_6.X a_8968_13760# VSS VSS sg13_lv_nmos ad=0.2886p pd=2.26u as=0.14875p ps=1.16u w=0.74u l=0.13u
x3087 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3088 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3089 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3090 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3091 a_16048_15454# sg13_inv_1_0.Y a_16108_15549# VDD sg13_lv_pmos ad=79.8f pd=0.8u as=0.204p ps=1.835u w=0.42u l=0.13u
x3092 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3093 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3094 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3095 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3096 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3097 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3098 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3099 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3100 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3101 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3102 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3103 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3104 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3105 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3106 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3107 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3108 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3109 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3110 a_13456_13942# a_13199_13799# a_13618_13722# VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=37.8f ps=0.6u w=0.42u l=0.13u
x3111 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3112 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3113 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3114 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3115 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3116 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3117 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3118 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3119 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3120 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3121 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3122 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3123 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3124 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3125 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3126 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3127 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3128 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3129 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3130 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3131 sg13_inv_1_1.Y sg13_inv_1_1.A VDD VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.3808p ps=2.92u w=1.12u l=0.13u
x3132 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3133 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3134 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3135 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3136 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3137 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3138 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3139 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3140 sg13_dfrbpq_1_3.Q a_16458_15532# VSS VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.1406p ps=1.12u w=0.74u l=0.13u
x3141 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3142 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3143 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3144 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3145 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3146 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3147 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3148 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3149 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3150 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3151 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3152 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3153 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3154 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3155 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3156 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3157 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3158 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3159 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3160 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3161 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3162 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3163 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3164 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3165 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3166 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3167 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3168 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3169 a_15599_16357# a_14757_16007# a_14340_16000# VDD sg13_lv_pmos ad=0.2048p pd=1.63u as=0.34p ps=2.68u w=1u l=0.13u
x3170 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3171 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3172 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3173 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3174 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3175 a_12650_15532# sg13_nor2_1_0.A VDD VDD sg13_lv_pmos ad=0.1176p pd=1.33u as=0.4032p ps=2.96u w=1.12u l=0.13u
x3176 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3177 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3178 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3179 a_14128_16966# a_13871_16823# a_14290_16746# VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=37.8f ps=0.6u w=0.42u l=0.13u
x3180 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3181 sg13_dfrbpq_1_6.D sg13_a22oi_1_0.B2 a_15096_17064# VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.15u
x3182 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3183 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3184 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3185 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3186 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3187 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3188 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3189 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3190 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3191 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3192 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3193 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3194 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3195 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3196 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3197 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3198 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3199 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3200 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3201 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3202 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3203 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3204 a_13871_16823# a_13029_16725# a_12612_17064# VDD sg13_lv_pmos ad=0.2048p pd=1.63u as=0.34p ps=2.68u w=1u l=0.13u
x3205 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3206 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3207 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3208 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3209 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3210 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3211 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3212 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3213 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3214 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3215 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3216 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3217 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3218 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3219 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3220 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3221 a_13401_14037# a_12459_13844# a_13199_13799# VDD sg13_lv_pmos ad=93.45f pd=0.865u as=0.2048p ps=1.63u w=0.42u l=0.13u
x3222 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3223 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3224 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3225 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3226 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3227 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3228 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3229 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3230 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3231 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3232 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3233 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3234 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3235 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3236 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3237 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3238 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3239 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3240 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3241 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3242 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3243 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3244 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3245 a_16294_14484# sg13_a21o_1_1.A2 VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0.19p ps=1.38u w=1u l=0.13u
x3246 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3247 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3248 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3249 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3250 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3251 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3252 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3253 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3254 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3255 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3256 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3257 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3258 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3259 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3260 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3261 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3262 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3263 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3264 VSS sg13_inv_2_1.A sg13_a21o_1_1.A2 VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.1406p ps=1.12u w=0.74u l=0.13u
x3265 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3266 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3267 VDD sg13_buf_1_4.A a_13768_10736# VDD sg13_lv_pmos ad=0.2114p pd=1.54u as=0.2856p ps=2.36u w=0.84u l=0.13u
x3268 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3269 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3270 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3271 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3272 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3273 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3274 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3275 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3276 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3277 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3278 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3279 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3280 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3281 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3282 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3283 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3284 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3285 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3286 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3287 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3288 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3289 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3290 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3291 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3292 a_13996_14607# a_13936_14726# a_13881_14607# VDD sg13_lv_pmos ad=0.204p pd=1.835u as=93.45f ps=0.865u w=0.42u l=0.13u
x3293 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3294 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3295 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3296 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3297 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3298 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3299 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3300 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3301 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3302 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3303 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3304 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3305 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3306 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3307 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3308 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3309 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3310 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3311 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3312 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3313 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3314 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3315 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3316 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3317 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3318 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3319 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3320 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3321 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3322 VDD adc_done a_17800_15272# VDD sg13_lv_pmos ad=0.2114p pd=1.54u as=0.2856p ps=2.36u w=0.84u l=0.13u
x3323 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3324 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3325 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3326 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3327 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3328 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3329 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3330 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3331 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3332 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3333 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3334 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3335 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3336 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3337 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3338 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3339 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3340 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3341 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3342 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3343 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3344 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3345 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3346 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3347 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3348 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3349 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3350 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3351 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3352 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3353 VDD sg13_inv_2_1.A a_16735_15972# VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2744p ps=1.61u w=1.12u l=0.13u
x3354 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3355 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3356 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3357 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3358 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3359 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3360 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3361 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3362 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3363 a_14340_15234# sg13_dfrbpq_1_3.D a_14246_15234# VSS sg13_lv_nmos ad=60.89999f pd=0.71u as=0.1428p ps=1.52u w=0.42u l=0.13u
x3364 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3365 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3366 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3367 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3368 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3369 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3370 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3371 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3372 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3373 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3374 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3375 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3376 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3377 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3378 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3379 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3380 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3381 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3382 VDD a_13459_12404# sg13_a21o_1_0.X VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.3808p ps=2.92u w=1.12u l=0.13u
x3383 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3384 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3385 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3386 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3387 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3388 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3389 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3390 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3391 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3392 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3393 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3394 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3395 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3396 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3397 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3398 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3399 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3400 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3401 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3402 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3403 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3404 a_14437_17878# sg13_a21oi_1_0.A1 VSS VSS sg13_lv_nmos ad=0.1406p pd=1.12u as=0.14505p ps=1.15u w=0.74u l=0.13u
x3405 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3406 a_14246_13722# sg13_and2_1_0.X VDD VDD sg13_lv_pmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
x3407 VSS sg13_inv_1_0.Y a_14340_13722# VSS sg13_lv_nmos ad=0.1626p pd=1.415u as=60.89999f ps=0.71u w=0.42u l=0.13u
x3408 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3409 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3410 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3411 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3412 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3413 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3414 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3415 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3416 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3417 a_15993_14037# a_15051_13844# a_15791_13799# VDD sg13_lv_pmos ad=93.45f pd=0.865u as=0.2048p ps=1.63u w=0.42u l=0.13u
x3418 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3419 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3420 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3421 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3422 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3423 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3424 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3425 a_11364_16421# a_11076_16000# a_11302_16421# VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=37.8f ps=0.6u w=0.42u l=0.13u
x3426 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3427 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3428 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3429 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3430 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3431 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3432 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3433 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3434 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3435 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3436 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3437 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3438 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3439 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3440 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3441 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3442 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3443 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3444 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3445 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3446 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3447 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3448 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3449 a_13459_12404# sg13_buf_1_0.A VSS VSS sg13_lv_nmos ad=0.1216p pd=1.02u as=0.15745p ps=1.175u w=0.64u l=0.13u
x3450 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3451 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3452 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3453 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3454 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3455 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3456 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3457 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3458 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3459 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3460 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3461 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3462 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3463 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3464 a_12837_14495# sg13_dfrbpq_1_0.CLK a_13297_14837# VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.31732p ps=1.805u w=0.74u l=0.13u
x3465 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3466 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3467 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3468 Timer_en a_13768_10736# VDD VDD sg13_lv_pmos ad=0.42p pd=2.99u as=0.2114p ps=1.54u w=1.12u l=0.13u
x3469 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3470 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3471 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3472 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3473 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3474 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3475 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3476 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3477 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3478 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3479 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3480 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3481 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3482 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3483 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3484 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3485 VDD sg13_inv_1_0.Y a_12134_14922# VDD sg13_lv_pmos ad=0.36237p pd=2.605u as=79.8f ps=0.8u w=0.42u l=0.13u
x3486 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3487 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3488 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3489 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3490 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3491 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3492 a_14054_16434# a_14859_16007# a_14314_15964# VDD sg13_lv_pmos ad=0.1428p pd=1.52u as=79.8f ps=0.8u w=0.42u l=0.13u
x3493 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3494 VDD sg13_inv_2_1.A sg13_a21o_1_1.A2 VDD sg13_lv_pmos ad=0.3864p pd=2.93u as=0.2128p ps=1.5u w=1.12u l=0.13u
x3495 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3496 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3497 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3498 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3499 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3500 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3501 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3502 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3503 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3504 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3505 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3506 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3507 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3508 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3509 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3510 sg13_buf_1_4.A a_13866_14020# VSS VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.1406p ps=1.12u w=0.74u l=0.13u
x3511 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3512 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3513 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3514 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3515 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3516 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3517 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3518 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3519 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3520 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3521 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3522 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3523 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3524 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3525 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3526 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3527 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3528 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3529 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3530 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3531 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3532 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3533 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3534 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3535 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3536 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3537 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3538 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3539 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3540 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3541 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3542 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3543 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3544 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3545 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3546 VDD a_15791_15311# a_16458_15532# VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.3864p ps=2.93u w=1.12u l=0.13u
x3547 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3548 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3549 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3550 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3551 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3552 a_11364_16421# a_11595_16007# a_11050_15964# VSS sg13_lv_nmos ad=0.2373p pd=1.97u as=79.8f ps=0.8u w=0.42u l=0.13u
x3553 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3554 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3555 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3556 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3557 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3558 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3559 a_10790_16434# sg13_dfrbpq_1_4.D VDD VDD sg13_lv_pmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
x3560 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3561 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3562 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3563 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3564 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3565 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3566 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3567 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3568 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3569 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3570 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3571 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3572 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3573 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3574 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3575 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3576 VDD sg13_inv_1_0.Y a_12326_16746# VDD sg13_lv_pmos ad=0.36237p pd=2.605u as=79.8f ps=0.8u w=0.42u l=0.13u
x3577 a_13881_14607# a_12939_14495# a_13679_14845# VDD sg13_lv_pmos ad=93.45f pd=0.865u as=0.2048p ps=1.63u w=0.42u l=0.13u
x3578 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3579 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3580 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3581 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3582 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3583 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3584 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3585 VDD sg13_o21ai_1_0.B1 sg13_dfrbpq_1_6.D VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.15u
x3586 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3587 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3588 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3589 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3590 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3591 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3592 a_14889_15625# a_14532_15552# VDD VDD sg13_lv_pmos ad=63f pd=0.72u as=0.1563p ps=1.22u w=0.42u l=0.13u
x3593 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3594 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3595 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3596 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3597 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3598 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3599 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3600 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3601 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3602 sc_en a_14440_5412# VDD VDD sg13_lv_pmos ad=0.42p pd=2.99u as=0.2114p ps=1.54u w=1.12u l=0.13u
x3603 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3604 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3605 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3606 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3607 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3608 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3609 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3610 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3611 VSS uart_busy a_15976_25068# VSS sg13_lv_nmos ad=0.14875p pd=1.16u as=0.187p ps=1.78u w=0.55u l=0.13u
x3612 a_11654_13722# sg13_a21o_1_0.X VDD VDD sg13_lv_pmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
x3613 sg13_a21oi_1_0.A2 a_13960_25068# VSS VSS sg13_lv_nmos ad=0.2886p pd=2.26u as=0.14875p ps=1.16u w=0.74u l=0.13u
x3614 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3615 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3616 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3617 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3618 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3619 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3620 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3621 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3622 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3623 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3624 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3625 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3626 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3627 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3628 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3629 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3630 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3631 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3632 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3633 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3634 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3635 VSS sg13_inv_1_0.Y a_14148_16434# VSS sg13_lv_nmos ad=0.1626p pd=1.415u as=60.89999f ps=0.71u w=0.42u l=0.13u
x3636 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3637 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3638 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3639 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3640 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3641 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3642 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3643 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3644 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3645 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3646 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3647 VSS wake_up_sg a_10024_15996# VSS sg13_lv_nmos ad=0.14875p pd=1.16u as=0.187p ps=1.78u w=0.55u l=0.13u
x3648 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3649 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3650 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3651 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3652 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3653 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3654 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3655 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3656 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3657 a_12708_14909# a_12939_14495# a_12394_14452# VSS sg13_lv_nmos ad=0.2373p pd=1.97u as=79.8f ps=0.8u w=0.42u l=0.13u
x3658 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3659 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3660 a_15096_17064# sg13_o21ai_1_0.A1 VDD VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.3808p ps=2.92u w=1.12u l=0.15u
x3661 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3662 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3663 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3664 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3665 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3666 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3667 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3668 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3669 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3670 sg13_nor2_1_0.A a_10024_15996# VSS VSS sg13_lv_nmos ad=0.2886p pd=2.26u as=0.14875p ps=1.16u w=0.74u l=0.13u
x3671 VSS sg13_inv_1_0.Y a_12420_16746# VSS sg13_lv_nmos ad=0.1626p pd=1.415u as=60.89999f ps=0.71u w=0.42u l=0.13u
x3672 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3673 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3674 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3675 VDD uart_done a_13960_25068# VDD sg13_lv_pmos ad=0.2114p pd=1.54u as=0.2856p ps=2.36u w=0.84u l=0.13u
x3676 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3677 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3678 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3679 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3680 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3681 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3682 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3683 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3684 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3685 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3686 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3687 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3688 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3689 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3690 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3691 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3692 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3693 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3694 a_13499_15996# sg13_a21oi_1_0.A2 VDD VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
x3695 sg13_dfrbpq_1_1.Q a_16458_14020# VSS VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.1406p ps=1.12u w=0.74u l=0.13u
x3696 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3697 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3698 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3699 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3700 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3701 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3702 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3703 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3704 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3705 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3706 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3707 VDD sg13_inv_1_0.Y a_11050_15964# VDD sg13_lv_pmos ad=0.1563p pd=1.22u as=0.147p ps=1.54u w=0.42u l=0.13u
x3708 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3709 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3710 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3711 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3712 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3713 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3714 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3715 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3716 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3717 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3718 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3719 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3720 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3721 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3722 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3723 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3724 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3725 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3726 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3727 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3728 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3729 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3730 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3731 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3732 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3733 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3734 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3735 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3736 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3737 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3738 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3739 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3740 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3741 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3742 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3743 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3744 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3745 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3746 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3747 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3748 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3749 sg13_nor2_1_0.B a_13002_15996# VSS VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.1406p ps=1.12u w=0.74u l=0.13u
x3750 sg13_o21ai_1_0.B1 sg13_a21oi_1_0.A1 VDD VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2198p ps=1.53u w=1.12u l=0.13u
x3751 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3752 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3753 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3754 clk_gating_en a_14632_4688# VSS VSS sg13_lv_nmos ad=0.2886p pd=2.26u as=0.14875p ps=1.16u w=0.74u l=0.13u
x3755 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3756 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3757 VDD sg13_inv_1_0.Y a_10790_16434# VDD sg13_lv_pmos ad=0.36237p pd=2.605u as=79.8f ps=0.8u w=0.42u l=0.13u
x3758 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3759 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3760 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3761 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3762 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3763 VDD sg13_inv_1_0.Y a_14246_15234# VDD sg13_lv_pmos ad=0.36237p pd=2.605u as=79.8f ps=0.8u w=0.42u l=0.13u
x3764 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3765 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3766 VSS VDD VSS VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
x3767 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3768 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3769 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3770 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3771 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3772 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3773 sg13_dfrbpq_1_4.D sg13_nor2_1_0.Y VSS VSS sg13_lv_nmos ad=0.1406p pd=1.12u as=0.2516p ps=2.16u w=0.74u l=0.13u
x3774 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3775 VDD a_16051_14746# sg13_dfrbpq_1_3.D VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.3808p ps=2.92u w=1.12u l=0.13u
x3776 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
x3777 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3778 VSS VDD VSS VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
x3779 VDD VSS VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
x3780 VSS a_15856_16238# a_15505_16357# VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
x3781 VDD VSS VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
C0 a_17006_16388# sg13_dfrbpq_1_5.Q 0
C1 a_14235_17564# sg13_o21ai_1_0.B1 0.29113f
C2 a_13960_4782# a_14144_4782# 0.0524f
C3 a_14889_15625# sg13_inv_1_1.A 0
C4 a_17024_13854# VDD 0.06319f
C5 a_15791_13799# a_16051_14746# 0
C6 a_12459_13844# VDD 0.19509f
C7 a_12134_14922# a_12777_14531# 0.00801f
C8 a_12837_14495# a_13679_14845# 0.00307f
C9 a_12708_14909# a_12939_14495# 0.12701f
C10 uart_en sg13_buf_1_0.A 0.03977f
C11 a_13866_14020# sg13_inv_1_0.Y 0.01461f
C12 a_13002_15996# sg13_inv_1_1.Y 0
C13 adc_done sg13_a21o_1_1.A2 0
C14 sg13_dfrbpq_1_5.Q a_15680_16878# 0.01758f
C15 a_15051_15356# a_16048_15454# 0.02979f
C16 sg13_buf_1_0.A a_13576_4688# 0.2758f
C17 sg13_dfrbpq_1_6.D a_13864_16426# 0.00193f
C18 a_12612_17064# sg13_nor2_1_0.Y 0.00461f
C19 a_14340_16000# a_15599_16357# 0.01529f
C20 a_14757_16007# a_15856_16238# 0
C21 a_15993_14037# sg13_dfrbpq_1_1.Q 0
C22 a_13105_13799# a_12459_13844# 0.00647f
C23 a_13866_14020# a_13199_13799# 0.0894f
C24 uart_done a_13960_25068# 0.26647f
C25 a_12650_15532# sg13_nor2_1_0.Y 0.01296f
C26 a_13516_14037# VDD 0.00769f
C27 a_12900_16759# sg13_nor2_1_0.Y 0.0025f
C28 a_13679_14845# a_14346_14484# 0.0894f
C29 a_13936_14726# a_13585_14845# 0.008f
C30 sg13_buf_1_0.A a_13960_4572# 0.00147f
C31 a_13499_15996# sg13_a21oi_1_0.A2 0.07879f
C32 sg13_a22oi_1_0.B2 sg13_inv_1_1.Y 0.0025f
C33 a_15051_15356# a_15409_15255# 0.00104f
C34 a_14949_15213# a_15697_15311# 0.01058f
C35 a_16048_15454# a_16108_15549# 0.01042f
C36 a_15791_15311# a_16458_15532# 0.0894f
C37 sg13_inv_1_1.A a_12612_17064# 0
C38 a_14340_16000# sg13_dfrbpq_1_4.D 0
C39 a_16832_15366# sg13_inv_1_1.A 0.00394f
C40 sg13_nor2_1_0.A a_11493_16007# 0.00154f
C41 a_17024_13644# sg13_dfrbpq_1_1.Q 0.00102f
C42 sg13_a21oi_1_0.A1 a_13029_16725# 0.00184f
C43 a_13585_14845# sg13_buf_1_0.A 0
C44 a_12650_15532# sg13_inv_1_1.A 0
C45 a_15496_16668# sg13_dfrbpq_1_6.D 0.00618f
C46 a_9728_13854# VDD 0.10036f
C47 a_15051_15356# sg13_dfrbpq_1_0.CLK 0.04384f
C48 a_13960_25068# a_13856_25154# 0.00624f
C49 a_14506_15457# sg13_a21oi_1_0.A1 0
C50 adc_done a_25856_16668# 0
C51 a_15791_15311# a_16210_15234# 0.00174f
C52 a_16048_15454# a_15697_15311# 0.008f
C53 sg13_o21ai_1_0.A1 a_15496_16668# 0.00237f
C54 a_16266_15996# sg13_dfrbpq_1_3.Q 0.01003f
C55 a_14144_17938# sg13_a21oi_1_0.A2 0.00228f
C56 sg13_a22oi_1_0.B2 a_15916_16119# 0.00187f
C57 a_13401_14037# sg13_a21o_1_0.X 0
C58 a_14144_17594# VDD 0.08419f
C59 a_12326_16746# a_13871_16823# 0
C60 sg13_inv_1_1.A sg13_dfrbpq_1_5.Q 0.11359f
C61 sg13_a22oi_1_0.B2 a_15680_16668# 0
C62 sg13_nor2_1_0.A a_12136_16878# 0
C63 a_14073_17061# a_13871_16823# 0.00689f
C64 a_16108_15549# sg13_dfrbpq_1_0.CLK 0.00139f
C65 a_14061_12256# sg13_inv_1_0.Y 0
C66 a_12754_16434# sg13_nor2_1_0.Y 0
C67 adc_start a_17696_15156# 0
C68 a_13459_12404# a_13702_12532# 0.13617f
C69 sg13_dfrbpq_1_4.D sg13_a21oi_1_0.A2 0.00432f
C70 a_11848_15366# sg13_nor2_1_0.A 0.03085f
C71 a_13864_16082# a_14054_16434# 0.00201f
C72 a_14054_16434# a_13679_14845# 0
C73 sg13_a21oi_1_0.A1 a_11953_16349# 0
C74 a_12394_14452# VDD 0.10067f
C75 a_12326_16746# a_13489_17042# 0
C76 a_12612_17064# a_13131_16868# 0.34114f
C77 wake_up_sg VDD 1.55825f
C78 a_15697_15311# sg13_dfrbpq_1_0.CLK 0.00441f
C79 sg13_nor2b_1_0.Y sg13_nor2_1_0.Y 0.00972f
C80 a_13489_16767# a_12612_17064# 0.01835f
C81 a_12900_16759# a_13131_16868# 0.12701f
C82 a_13472_4572# VDD 0
C83 a_16430_14832# VDD 0
C84 sg13_dfrbpq_1_3.D a_16832_15366# 0
C85 a_14532_15552# sg13_o21ai_1_0.A1 0
C86 uart_busy tx_start 0.13424f
C87 a_13499_15996# VDD 0.26397f
C88 a_12900_16759# a_13489_16767# 0
C89 a_13936_14726# VDD 0.17826f
C90 sg13_dfrbpq_1_1.Q a_16832_15156# 0
C91 sg13_a22oi_1_0.B2 a_15505_16357# 0.00763f
C92 a_14949_15213# sg13_inv_2_1.A 0
C93 sg13_a22oi_1_0.B2 tx_start 0.05338f
C94 a_14949_15213# sg13_a22oi_1_0.B2 0.00126f
C95 a_14144_17938# VDD 0.00264f
C96 a_13192_12342# sg13_a21o_1_0.X 0.03677f
C97 a_15791_15311# sg13_o21ai_1_0.A1 0
C98 a_15599_16357# VDD 0.18329f
C99 sg13_dfrbpq_1_3.D a_14246_13722# 0.00156f
C100 sg13_dfrbpq_1_3.D sg13_dfrbpq_1_5.Q 0
C101 sg13_dfrbpq_1_0.CLK a_11493_16007# 0.27541f
C102 a_15217_15998# sg13_inv_1_0.Y 0.01659f
C103 sg13_buf_1_0.A VDD 2.76775f
C104 sg13_dfrbpq_1_6.D a_13871_16823# 0.02117f
C105 a_16048_15454# sg13_inv_2_1.A 0.00118f
C106 sg13_dfrbpq_1_1.Q a_16294_14484# 0.08523f
C107 sg13_o21ai_1_0.A1 a_13871_16823# 0
C108 a_14538_17044# a_14128_16966# 0.10373f
C109 a_14889_14113# sg13_dfrbpq_1_0.CLK 0
C110 a_16048_15454# sg13_a22oi_1_0.B2 0
C111 a_13105_13799# sg13_buf_1_0.A 0.00141f
C112 a_14889_15625# sg13_inv_1_0.Y 0
C113 a_13864_16082# sg13_inv_1_1.Y 0.04058f
C114 a_14061_12256# timer_done 0
C115 a_12326_16746# sg13_nor2_1_0.B 0
C116 sg13_dfrbpq_1_4.D VDD 0.42835f
C117 sg13_nor2_1_0.A a_11914_13945# 0
C118 a_14246_13722# a_14949_13701# 0.02454f
C119 sg13_dfrbpq_1_0.CLK a_13002_15996# 0.01183f
C120 a_11076_16000# a_11493_16007# 0.37384f
C121 sg13_inv_1_1.Y a_13679_14845# 0
C122 sg13_dfrbpq_1_6.D a_13489_17042# 0.00234f
C123 a_12136_16878# sg13_dfrbpq_1_0.CLK 0.00266f
C124 a_14340_16000# a_15680_16878# 0
C125 a_14757_16007# a_15496_16878# 0.00238f
C126 a_17128_13760# sg13_dfrbpq_1_0.CLK 0
C127 a_13777_16823# sg13_dfrbpq_1_6.D 0.00577f
C128 a_14538_17044# sg13_dfrbpq_1_0.CLK 0
C129 a_13601_16344# sg13_a21oi_1_0.A2 0.00205f
C130 a_14532_14040# a_15791_13799# 0.01529f
C131 sg13_dfrbpq_1_3.Q sg13_dfrbpq_1_1.Q 0.15484f
C132 sg13_buf_1_5.X Timer_en 0.02836f
C133 a_11848_15366# sg13_dfrbpq_1_0.CLK 0
C134 a_11364_16421# a_11595_16007# 0.12701f
C135 a_11493_16007# a_12335_16357# 0.00307f
C136 sg13_dfrbpq_1_3.D a_14820_13735# 0
C137 a_10790_16434# a_11433_16043# 0.00801f
C138 a_14538_17044# a_14290_16746# 0
C139 sg13_inv_2_1.A sg13_dfrbpq_1_0.CLK 0.0041f
C140 a_12136_16878# a_11076_16000# 0
C141 sg13_a22oi_1_0.B2 sg13_dfrbpq_1_0.CLK 0.22482f
C142 sg13_inv_1_0.Y a_12612_17064# 0.40714f
C143 a_12586_16969# a_13029_16725# 0.02242f
C144 sg13_dfrbpq_1_0.CLK a_12817_14018# 0.00251f
C145 sg13_nor2_1_0.A a_12420_14488# 0
C146 a_12046_15276# a_11493_16007# 0.00159f
C147 a_11848_15366# a_11076_16000# 0
C148 a_12900_16759# sg13_inv_1_0.Y 0.00396f
C149 a_15051_13844# a_15993_14037# 0
C150 a_14532_14040# a_14758_13735# 0.0052f
C151 a_14949_13701# a_14820_13735# 0.01562f
C152 a_12335_16357# a_13002_15996# 0.0894f
C153 a_12592_16238# a_12241_16357# 0.008f
C154 a_12650_15532# sg13_inv_1_0.Y 0.00356f
C155 timer_done sc_en 0.27424f
C156 sg13_dfrbpq_1_3.Q a_15801_16119# 0
C157 sg13_dfrbpq_1_6.D a_12592_16238# 0.0019f
C158 sc_en a_14632_4688# 0.04835f
C159 sg13_inv_1_1.A a_17696_15366# 0
C160 a_12228_13735# VDD 0.00693f
C161 sg13_nor2b_1_0.Y a_11595_16007# 0.00132f
C162 a_13864_16426# a_14054_16434# 0.00404f
C163 sg13_dfrbpq_1_5.Q sg13_inv_1_0.Y 0.00147f
C164 a_12241_16357# sg13_nor2_1_0.B 0
C165 a_16458_14020# a_17128_13760# 0
C166 a_14246_13722# sg13_inv_1_0.Y 0.11428f
C167 sg13_a21o_1_0.A2 sg13_buf_1_5.X 0.29471f
C168 a_12046_15276# a_12136_16878# 0
C169 sg13_and2_1_0.X a_14949_13701# 0.00142f
C170 a_14506_13945# a_15051_13844# 0.01f
C171 a_14340_16000# sg13_inv_1_1.A 0.00147f
C172 sg13_dfrbpq_1_6.D sg13_nor2_1_0.B 0.00235f
C173 sg13_inv_1_0.Y a_11364_16421# 0
C174 a_12046_15276# a_11848_15366# 0.01393f
C175 sg13_a21oi_1_0.A1 a_14757_16007# 0.00668f
C176 sg13_o21ai_1_0.B1 a_13871_16823# 0.00207f
C177 a_13480_10830# sg13_buf_1_0.A 0.00926f
C178 a_14340_13722# sg13_inv_1_0.Y 0
C179 a_15784_14570# VDD 0.16488f
C180 a_14820_13735# a_15409_13743# 0
C181 sg13_and2_1_0.X a_16048_13942# 0
C182 a_17024_13854# a_17128_13760# 0.00624f
C183 a_13601_16344# VDD 0
C184 a_13618_13722# a_13456_13942# 0.00188f
C185 a_15599_16357# a_16018_16434# 0.00174f
C186 a_14859_16007# a_15217_15998# 0.02138f
C187 a_13881_14607# VDD 0.00138f
C188 sg13_inv_1_0.Y a_12754_16434# 0.00114f
C189 sg13_a21oi_1_0.A1 a_15217_16349# 0
C190 sg13_a21oi_1_0.A1 a_14144_23642# 0.02298f
C191 a_15791_15311# a_16294_14484# 0
C192 sg13_nor2b_1_0.Y a_11940_14040# 0
C193 a_14152_5498# sg13_buf_1_0.A 0.01194f
C194 tx_start a_13960_25068# 0.00332f
C195 a_14532_15552# sg13_dfrbpq_1_3.Q 0
C196 a_15051_15356# a_15599_16357# 0
C197 a_14820_13735# sg13_inv_1_0.Y 0.00158f
C198 sg13_nor2b_1_0.Y sg13_inv_1_0.Y 0.18535f
C199 a_17006_16388# VDD 0
C200 sg13_and2_1_0.X a_15409_13743# 0
C201 sg13_buf_1_5.X sg13_a21o_1_0.X 0
C202 a_14061_12256# a_13866_14020# 0
C203 a_12459_13844# a_12817_14018# 0.02138f
C204 a_11654_13722# a_11748_13722# 0.00716f
C205 a_13702_12532# VDD 0.34097f
C206 a_15680_16878# VDD 0.07064f
C207 sg13_dfrbpq_1_0.CLK a_12420_14488# 0.10683f
C208 a_16840_13854# sg13_dfrbpq_1_0.CLK 0
C209 sg13_a21o_1_1.A2 a_16051_14746# 0.00145f
C210 a_15791_15311# sg13_dfrbpq_1_3.Q 0.00902f
C211 sg13_and2_1_0.X sg13_inv_1_0.Y 0.17346f
C212 sg13_dfrbpq_1_3.D a_14340_16000# 0
C213 a_13459_12404# sg13_inv_1_0.Y 0.00131f
C214 sg13_inv_1_0.Y a_11464_13644# 0.00247f
C215 sg13_inv_1_1.Y a_13996_14607# 0
C216 a_13459_12404# a_13199_13799# 0
C217 a_13864_16082# sg13_dfrbpq_1_0.CLK 0.01121f
C218 a_25856_11546# VDD 0.0583f
C219 sg13_dfrbpq_1_0.CLK a_13679_14845# 0.0105f
C220 a_10024_15996# VDD 0.26883f
C221 wake_up_sg a_11493_16007# 0
C222 sg13_nor2_1_0.Y VDD 0.44431f
C223 sg13_a21oi_1_0.A1 a_14314_15964# 0.00473f
C224 a_13131_16868# sg13_a21oi_1_0.A2 0.03088f
C225 a_11914_13945# a_12459_13844# 0.01f
C226 sg13_a21o_1_0.X a_11654_13722# 0.27608f
C227 a_14152_5842# VDD 0.00916f
C228 a_16266_15996# sg13_dfrbpq_1_0.CLK 0.00152f
C229 Timer_en a_14248_4688# 0.00655f
C230 a_12592_16238# a_12837_14495# 0
C231 a_12335_16357# a_12420_14488# 0
C232 reset VDD 1.34688f
C233 a_14859_16007# sg13_dfrbpq_1_5.Q 0
C234 a_14246_15234# VDD 0.79999f
C235 a_14336_5498# VDD 0.06961f
C236 a_16840_13854# a_16458_14020# 0.01012f
C237 a_13871_16823# a_14054_16434# 0
C238 sg13_nor2b_1_0.Y a_12134_14922# 0.27178f
C239 sg13_inv_1_0.Y a_11464_13854# 0.01456f
C240 sg13_inv_1_1.A VDD 0.53573f
C241 sg13_a21o_1_0.A2 sg13_a21o_1_0.X 0
C242 sg13_a21o_1_0.X a_11748_13722# 0
C243 sg13_nor2_1_0.B a_12837_14495# 0.0021f
C244 Timer_en a_14144_4572# 0.00131f
C245 a_14340_15234# VDD 0
C246 a_12459_13844# a_12420_14488# 0
C247 a_12357_13701# a_12837_14495# 0.00173f
C248 a_16840_13854# a_17024_13854# 0.0524f
C249 a_12420_16746# VDD 0
C250 sg13_dfrbpq_1_4.D a_11493_16007# 0.0131f
C251 a_16735_16388# sg13_a21o_1_1.A2 0
C252 a_15051_15356# a_15784_14570# 0
C253 a_14820_15247# VDD 0.00858f
C254 a_14340_16000# sg13_inv_1_0.Y 0.38254f
C255 a_14532_15552# sg13_inv_1_1.Y 0
C256 a_14506_15457# a_14314_15964# 0
C257 a_15856_16238# sg13_o21ai_1_0.A1 0
C258 sg13_inv_1_0.Y a_12646_14909# 0
C259 a_13456_13942# a_12837_14495# 0
C260 sg13_dfrbpq_1_4.D a_13002_15996# 0.01012f
C261 a_13131_16868# VDD 0.19128f
C262 a_12136_16878# sg13_dfrbpq_1_4.D 0
C263 sg13_a22oi_1_0.B2 a_15599_16357# 0.02317f
C264 a_16048_15454# sg13_dfrbpq_1_1.Q 0.00107f
C265 a_14628_16421# sg13_inv_1_0.Y 0.00138f
C266 sg13_dfrbpq_1_3.D VDD 0.48775f
C267 a_13489_16767# VDD 0
C268 a_13768_10736# a_14152_10736# 0.0015f
C269 sg13_a21oi_1_0.A1 a_14998_16742# 0.02723f
C270 sg13_inv_1_0.Y a_13585_14845# 0.00211f
C271 a_11848_15366# sg13_dfrbpq_1_4.D 0.0021f
C272 clk sg13_dfrbpq_1_0.CLK 0.06214f
C273 sg13_inv_1_1.A a_16735_15972# 0.1784f
C274 a_13199_13799# a_13585_14845# 0
C275 a_10884_16434# VDD 0
C276 a_13871_16823# sg13_inv_1_1.Y 0.001f
C277 a_13866_14020# a_14246_13722# 0
C278 sg13_inv_1_0.Y sg13_a21oi_1_0.A2 0.02943f
C279 a_15697_15311# a_15784_14570# 0
C280 a_14949_13701# VDD 0.2642f
C281 Timer_en adc_en 1.57613f
C282 a_11595_16007# VDD 0.18782f
C283 timer_done uart_en 0.76759f
C284 sg13_dfrbpq_1_0.CLK sg13_dfrbpq_1_1.Q 0.03476f
C285 sg13_buf_1_5.X sg13_buf_1_4.A 0.45745f
C286 timer_done a_13576_4688# 0
C287 uart_en a_14632_4688# 0.08855f
C288 a_16048_13942# VDD 0.16276f
C289 a_13777_16823# sg13_inv_1_1.Y 0.00102f
C290 sg13_dfrbpq_1_0.CLK a_13996_14607# 0.00143f
C291 a_14336_5842# a_14440_5412# 0
C292 sg13_dfrbpq_1_5.Q a_15784_14914# 0
C293 a_12394_14452# a_12420_14488# 0.36952f
C294 a_16210_13722# a_15697_13799# 0
C295 a_11953_15998# VDD 0.00645f
C296 a_11914_13945# sg13_buf_1_0.A 0
C297 a_15801_16119# sg13_dfrbpq_1_0.CLK 0.00134f
C298 Timer_en sg13_buf_1_4.A 0.00486f
C299 a_14152_5498# a_14336_5498# 0.0524f
C300 a_14532_15552# a_14949_15213# 0.3749f
C301 a_14246_15234# a_15051_15356# 0.097f
C302 timer_done a_13960_4572# 0
C303 a_15409_13743# VDD 0.00143f
C304 a_15051_15356# sg13_inv_1_1.A 0.02272f
C305 a_14248_4688# a_14144_4572# 0
C306 a_14235_17564# a_14144_17594# 0.00761f
C307 a_13192_12132# sg13_dfrbpq_1_0.CLK 0
C308 a_12837_14495# a_12939_14495# 0.47795f
C309 a_12420_14488# a_13936_14726# 0.00139f
C310 a_15496_16668# sg13_dfrbpq_1_0.CLK 0.00118f
C311 a_11940_14040# VDD 0.08626f
C312 a_15688_25154# VDD 0.1353f
C313 a_17024_13644# adc_start 0
C314 a_15791_13799# sg13_a21o_1_1.A2 0.00194f
C315 a_14246_15234# a_16108_15549# 0
C316 a_14532_15552# a_16048_15454# 0.00242f
C317 a_14949_15213# a_15791_15311# 0.00332f
C318 a_13105_13799# a_11940_14040# 0.43239f
C319 a_12817_13743# a_12357_13701# 0.02396f
C320 sg13_inv_1_0.Y VDD 10.0839f
C321 a_13866_14020# sg13_and2_1_0.X 0.01133f
C322 a_14340_16000# a_14859_16007# 0.34102f
C323 a_14757_16007# a_15217_16349# 0.02396f
C324 a_13499_15996# a_13864_16082# 0.01004f
C325 a_16458_14020# sg13_dfrbpq_1_1.Q 0.12431f
C326 a_9920_16082# sg13_dfrbpq_1_0.CLK 0.00209f
C327 a_16108_15549# sg13_inv_1_1.A 0.0031f
C328 a_13864_16082# a_13936_14726# 0
C329 a_13199_13799# VDD 0.18663f
C330 a_12420_14488# sg13_buf_1_0.A 0
C331 a_12837_14495# a_13297_14486# 0.01483f
C332 a_13936_14726# a_13679_14845# 0.34468f
C333 sg13_nor2_1_0.B sg13_inv_1_1.Y 0
C334 a_13105_13799# sg13_inv_1_0.Y 0.00532f
C335 sg13_a22oi_1_0.B2 a_15784_14570# 0
C336 sg13_buf_1_0.A a_13960_4782# 0.01025f
C337 sg13_a21o_1_0.A2 sg13_buf_1_4.A 0.5612f
C338 a_15791_15311# a_16048_15454# 0.34468f
C339 a_14532_15552# a_15409_15255# 0.01835f
C340 a_15051_15356# a_14820_15247# 0.12701f
C341 a_14628_16421# a_14859_16007# 0.12701f
C342 a_13105_13799# a_13199_13799# 0.28931f
C343 a_17024_13854# sg13_dfrbpq_1_1.Q 0.02574f
C344 sg13_dfrbpq_1_4.D a_12420_14488# 0
C345 a_15697_15311# sg13_inv_1_1.A 0
C346 sg13_nor2_1_0.A a_11050_15964# 0
C347 sg13_dfrbpq_1_3.D a_16018_16434# 0
C348 a_13679_14845# sg13_buf_1_0.A 0.00209f
C349 a_15496_16878# sg13_dfrbpq_1_6.D 0.02067f
C350 sg13_a21oi_1_0.A1 a_14073_17061# 0
C351 a_14532_15552# sg13_dfrbpq_1_0.CLK 0.09602f
C352 a_8776_13854# VDD 0.14617f
C353 a_11493_16007# sg13_nor2_1_0.Y 0
C354 a_14859_16007# sg13_a21oi_1_0.A2 0
C355 sg13_o21ai_1_0.A1 a_15496_16878# 0.00903f
C356 sg13_inv_2_1.A a_17006_16388# 0.00108f
C357 a_15856_16238# sg13_dfrbpq_1_3.Q 0.00142f
C358 a_15599_16357# a_16266_15996# 0.0894f
C359 sg13_dfrbpq_1_3.D a_15051_15356# 0.01234f
C360 a_13871_16823# a_14128_16966# 0.34468f
C361 a_13864_16082# sg13_dfrbpq_1_4.D 0.00113f
C362 a_12326_16746# a_12136_16668# 0.00404f
C363 a_14144_17938# a_14235_17564# 0
C364 a_12228_13735# a_11914_13945# 0.00463f
C365 sg13_nor2_1_0.A a_12592_16238# 0.00154f
C366 sg13_a21oi_1_0.A1 a_15096_17064# 0.00199f
C367 a_15791_15311# sg13_dfrbpq_1_0.CLK 0.00684f
C368 sg13_a22oi_1_0.B2 a_15680_16878# 0
C369 a_13459_12404# a_14061_12256# 0.00483f
C370 a_13002_15996# sg13_nor2_1_0.Y 0.05764f
C371 a_14061_12256# sg13_and2_1_0.X 0.10477f
C372 a_14757_16007# a_14314_15964# 0.02242f
C373 a_14949_15213# a_15051_13844# 0
C374 adc_en a_14248_4688# 0.02572f
C375 sg13_buf_1_4.A sg13_a21o_1_0.X 0
C376 sg13_dfrbpq_1_0.CLK a_13871_16823# 0
C377 sg13_nor2_1_0.A sg13_nor2_1_0.B 0.30504f
C378 a_12134_14922# VDD 0.79005f
C379 a_12326_16746# a_13029_16725# 0.02454f
C380 timer_done VDD 1.80756f
C381 a_14758_15247# sg13_dfrbpq_1_0.CLK 0
C382 a_14290_16746# a_13871_16823# 0.00174f
C383 a_13777_16823# a_14128_16966# 0.008f
C384 a_12900_16759# a_12612_17064# 0.43707f
C385 a_14632_4688# VDD 0.22656f
C386 sg13_nor2_1_0.A a_12357_13701# 0
C387 sg13_dfrbpq_1_3.D a_15697_15311# 0.02337f
C388 clk wake_up_sg 0.66497f
C389 sg13_a21oi_1_0.A1 a_12241_16357# 0
C390 a_12537_16119# VDD 0
C391 adc_en a_14144_4572# 0
C392 a_13489_17042# sg13_dfrbpq_1_0.CLK 0.00171f
C393 sg13_a21oi_1_0.A1 sg13_dfrbpq_1_6.D 0.15291f
C394 a_13297_14837# VDD 0.00223f
C395 a_14246_15234# sg13_a22oi_1_0.B2 0
C396 sg13_buf_1_6.X VDD 0.42191f
C397 a_25768_4782# VDD 0.13597f
C398 sg13_a21oi_1_0.A1 sg13_o21ai_1_0.A1 0.05349f
C399 sg13_a21o_1_1.A2 a_17696_15156# 0
C400 a_15791_15311# a_16458_14020# 0
C401 a_16458_15532# a_15791_13799# 0
C402 a_15697_15311# a_14949_13701# 0
C403 sg13_inv_2_1.A sg13_inv_1_1.A 0.69879f
C404 a_16832_15366# sg13_dfrbpq_1_5.Q 0.00116f
C405 a_14859_16007# VDD 0.19257f
C406 a_13777_16823# a_14290_16746# 0
C407 a_12777_14531# VDD 0
C408 a_25768_23986# VDD 0.00121f
C409 sg13_a22oi_1_0.B2 sg13_inv_1_1.A 0.27599f
C410 sg13_dfrbpq_1_0.CLK a_11050_15964# 0.0126f
C411 tx_start a_15872_25154# 0
C412 sg13_dfrbpq_1_6.D a_12136_16668# 0.00154f
C413 sg13_dfrbpq_1_1.Q a_16430_14832# 0
C414 a_15051_13844# sg13_dfrbpq_1_0.CLK 0.03561f
C415 a_15496_16878# sg13_o21ai_1_0.B1 0.01551f
C416 a_14188_17061# a_13871_16823# 0.00247f
C417 a_15697_15311# a_16048_13942# 0
C418 a_15051_15356# sg13_inv_1_0.Y 0.4257f
C419 a_11050_15964# a_11076_16000# 0.36952f
C420 a_16294_14484# a_16051_14746# 0.13617f
C421 sg13_dfrbpq_1_3.D a_14889_14113# 0
C422 sg13_dfrbpq_1_0.CLK a_12592_16238# 0.0107f
C423 sg13_dfrbpq_1_6.D a_13029_16725# 0.01883f
C424 a_13679_14845# a_13881_14607# 0.00689f
C425 a_13936_14726# a_13996_14607# 0.01042f
C426 a_16108_14037# sg13_dfrbpq_1_0.CLK 0.00139f
C427 a_14757_16007# a_14998_16742# 0.00108f
C428 a_12838_16759# sg13_dfrbpq_1_6.D 0
C429 sg13_o21ai_1_0.A1 a_13029_16725# 0
C430 a_14820_15247# sg13_a22oi_1_0.B2 0
C431 a_16108_15549# sg13_inv_1_0.Y 0.01227f
C432 a_15599_16357# sg13_dfrbpq_1_1.Q 0
C433 a_15051_13844# a_15409_14018# 0.02138f
C434 a_14246_13722# a_14340_13722# 0.00716f
C435 a_11076_16000# a_12592_16238# 0.00139f
C436 a_11493_16007# a_11595_16007# 0.47795f
C437 a_14506_15457# sg13_o21ai_1_0.A1 0
C438 sg13_dfrbpq_1_0.CLK sg13_nor2_1_0.B 0.13788f
C439 sg13_nor2b_1_0.Y a_12650_15532# 0
C440 sg13_dfrbpq_1_3.Q a_16051_14746# 0.01675f
C441 sg13_buf_1_0.A a_13996_14607# 0.00194f
C442 a_12586_16969# a_12326_16746# 0.75507f
C443 sg13_nor2_1_0.A a_12228_14922# 0
C444 sg13_dfrbpq_1_3.D sg13_inv_2_1.A 0.00235f
C445 a_15697_15311# sg13_inv_1_0.Y 0
C446 sg13_dfrbpq_1_3.D sg13_a22oi_1_0.B2 0
C447 sg13_dfrbpq_1_0.CLK a_12357_13701# 0.27179f
C448 sc_en uart_en 1.13309f
C449 a_15599_16357# a_15801_16119# 0.00689f
C450 a_15856_16238# a_15916_16119# 0.01042f
C451 a_12592_16238# a_12335_16357# 0.34468f
C452 wake_up_sg a_9920_16082# 0.02391f
C453 a_11493_16007# a_11953_15998# 0.01483f
C454 a_11076_16000# sg13_nor2_1_0.B 0
C455 a_14246_13722# a_14820_13735# 0.31978f
C456 a_16210_13722# adc_start 0
C457 a_12136_16878# a_11595_16007# 0
C458 sg13_nor2_1_0.Y a_12420_14488# 0
C459 sg13_a21oi_1_0.A1 sg13_o21ai_1_0.B1 0.15249f
C460 a_13866_14020# VDD 0.38905f
C461 a_13192_12132# sg13_buf_1_0.A 0.00234f
C462 a_11848_15366# a_11595_16007# 0
C463 a_15791_13799# a_15993_14037# 0.00689f
C464 a_14152_5498# timer_done 0.00315f
C465 sg13_dfrbpq_1_0.CLK a_13456_13942# 0.01698f
C466 a_12335_16357# sg13_nor2_1_0.B 0.0028f
C467 a_14506_13945# a_14532_14040# 0.36952f
C468 sg13_and2_1_0.X a_14246_13722# 0.27646f
C469 a_14340_16000# a_15217_15998# 0
C470 a_12228_13735# a_12166_13735# 0
C471 sg13_inv_1_0.Y a_11493_16007# 0.04385f
C472 sg13_a21oi_1_0.A1 a_12837_14495# 0
C473 a_13768_10736# sg13_buf_1_0.A 0.04455f
C474 a_12046_15276# sg13_nor2_1_0.B 0.06176f
C475 a_14889_14113# sg13_inv_1_0.Y 0
C476 a_14246_15234# a_13679_14845# 0
C477 a_17800_15272# a_17696_15366# 0.00624f
C478 sg13_and2_1_0.X a_14340_13722# 0
C479 a_15856_16238# a_15505_16357# 0.008f
C480 a_15784_14914# VDD 0.00332f
C481 sg13_inv_1_0.Y a_13002_15996# 0.0033f
C482 sg13_inv_1_1.A a_13679_14845# 0.0016f
C483 sg13_a21oi_1_0.A1 a_14566_16421# 0
C484 uart_busy a_15688_25154# 0.00537f
C485 a_9920_16082# sg13_dfrbpq_1_4.D 0
C486 a_14336_5842# sg13_buf_1_0.A 0
C487 sg13_inv_1_0.Y a_12136_16878# 0.00135f
C488 a_12586_16969# sg13_dfrbpq_1_6.D 0.01319f
C489 sg13_nor2_1_0.B a_12459_13844# 0.00155f
C490 a_15051_15356# a_14859_16007# 0
C491 a_15688_25498# a_15976_25068# 0
C492 sg13_and2_1_0.X a_14820_13735# 0.00326f
C493 a_14532_15552# sg13_buf_1_0.A 0
C494 a_11848_15366# sg13_inv_1_0.Y 0.00334f
C495 a_14538_17044# sg13_inv_1_0.Y 0.00345f
C496 sg13_a22oi_1_0.B2 a_15688_25154# 0
C497 sg13_dfrbpq_1_3.Q a_16735_16388# 0.01722f
C498 a_16266_15996# sg13_inv_1_1.A 0.0029f
C499 a_14248_23556# sg13_a21oi_1_0.A2 0.00763f
C500 sg13_inv_2_1.A sg13_inv_1_0.Y 0
C501 a_11940_14040# a_12817_14018# 0
C502 a_11654_13722# a_12297_14113# 0.00801f
C503 a_12357_13701# a_12459_13844# 0.47622f
C504 sg13_a22oi_1_0.B2 sg13_inv_1_0.Y 0.01117f
C505 a_14912_16668# VDD 0
C506 a_14061_12256# VDD 0.41908f
C507 a_16048_15454# a_15856_16238# 0
C508 a_15791_15311# a_15599_16357# 0.00198f
C509 a_15784_14570# sg13_dfrbpq_1_1.Q 0.00226f
C510 sg13_inv_1_0.Y a_12817_14018# 0.02121f
C511 a_12969_17137# sg13_a21oi_1_0.A2 0
C512 a_12459_13844# a_13456_13942# 0.02979f
C513 a_12652_16119# sg13_dfrbpq_1_0.CLK 0
C514 a_13864_16082# a_13131_16868# 0
C515 a_7816_15996# VDD 0.31209f
C516 a_25856_11890# VDD 0
C517 a_11493_16007# a_12134_14922# 0
C518 wake_up_sg a_11050_15964# 0
C519 sg13_dfrbpq_1_0.CLK a_12939_14495# 0.04495f
C520 a_14340_16000# sg13_dfrbpq_1_5.Q 0.00102f
C521 a_14697_16043# a_14314_15964# 0.00333f
C522 sg13_a21oi_1_0.A1 a_14054_16434# 0.01545f
C523 sg13_dfrbpq_1_3.D a_13679_14845# 0.0039f
C524 a_12612_17064# sg13_a21oi_1_0.A2 0.05704f
C525 a_13456_13942# a_13516_14037# 0.01042f
C526 a_15856_16238# sg13_dfrbpq_1_0.CLK 0.00322f
C527 a_13480_10620# VDD 0.0024f
C528 sg13_dfrbpq_1_0.CLK a_13297_14486# 0.00692f
C529 a_12592_16238# a_12394_14452# 0
C530 a_12900_16759# sg13_a21oi_1_0.A2 0
C531 a_11914_13945# a_11940_14040# 0.36952f
C532 sc_en VDD 0.33721f
C533 a_14532_14040# a_14346_14484# 0
C534 sg13_inv_1_0.Y a_11914_13945# 0.26965f
C535 a_15217_15998# VDD 0.0078f
C536 a_13664_10830# sg13_buf_1_4.A 0.0219f
C537 a_12652_16119# a_12335_16357# 0.00247f
C538 a_14248_23556# VDD 0.28393f
C539 Timer_en a_14144_4782# 0.00275f
C540 a_15791_13799# a_16294_14484# 0
C541 sg13_nor2_1_0.B a_12394_14452# 0.0039f
C542 a_14757_16007# sg13_dfrbpq_1_6.D 0.00214f
C543 a_14889_15625# VDD 0
C544 a_14061_12256# a_14155_12256# 0.00273f
C545 a_14757_16007# sg13_o21ai_1_0.A1 0.00431f
C546 a_13499_15996# sg13_nor2_1_0.B 0
C547 sg13_dfrbpq_1_4.D a_11050_15964# 0.01923f
C548 a_12969_17137# VDD 0
C549 a_15217_16349# sg13_dfrbpq_1_6.D 0.00171f
C550 sg13_dfrbpq_1_3.Q a_15791_13799# 0.00135f
C551 a_14506_15457# a_14054_16434# 0
C552 a_14532_15552# a_15784_14570# 0
C553 a_17800_15272# VDD 0.26811f
C554 sg13_inv_1_0.Y a_12420_14488# 0.43912f
C555 sg13_inv_1_1.A sg13_dfrbpq_1_1.Q 0.02284f
C556 a_13199_13799# a_12420_14488# 0
C557 sg13_a21oi_1_0.A1 sg13_inv_1_1.Y 0.01806f
C558 sg13_dfrbpq_1_4.D a_12592_16238# 0.00649f
C559 a_12459_13844# a_12939_14495# 0
C560 sg13_inv_1_1.A a_13996_14607# 0
C561 a_12612_17064# VDD 0.07873f
C562 sg13_a22oi_1_0.B2 a_14859_16007# 0.02629f
C563 a_15791_15311# a_15784_14570# 0
C564 a_16832_15366# VDD 0.0815f
C565 a_13864_16082# sg13_inv_1_0.Y 0
C566 a_15505_16357# a_15496_16878# 0
C567 a_12900_16759# VDD 0.00678f
C568 sg13_inv_1_0.Y a_13679_14845# 0.14653f
C569 a_12650_15532# VDD 0.00804f
C570 a_13401_14037# sg13_dfrbpq_1_0.CLK 0.00344f
C571 a_16048_15454# a_16051_14746# 0.00142f
C572 a_10024_15996# a_9920_16082# 0.00624f
C573 sg13_inv_1_1.A a_15801_16119# 0
C574 a_12357_13701# sg13_buf_1_0.A 0
C575 a_13199_13799# a_13679_14845# 0
C576 a_16458_15532# sg13_a21o_1_1.A2 0.00151f
C577 sg13_dfrbpq_1_4.D sg13_nor2_1_0.B 0.15506f
C578 a_16266_15996# sg13_inv_1_0.Y 0
C579 a_14235_17564# sg13_inv_1_0.Y 0
C580 a_14246_13722# VDD 0.80131f
C581 sg13_dfrbpq_1_5.Q VDD 0.57264f
C582 a_16210_15234# sg13_a21o_1_1.A2 0
C583 a_13456_13942# sg13_buf_1_0.A 0.00985f
C584 a_16210_13722# a_15791_13799# 0.00174f
C585 a_11364_16421# VDD 0.00601f
C586 sg13_dfrbpq_1_6.D a_14314_15964# 0
C587 sg13_dfrbpq_1_3.D sg13_dfrbpq_1_1.Q 0.00524f
C588 sg13_dfrbpq_1_0.CLK a_16051_14746# 0.00338f
C589 a_14757_16007# sg13_o21ai_1_0.B1 0
C590 a_14506_15457# sg13_inv_1_1.Y 0
C591 a_14340_13722# VDD 0
C592 a_12134_14922# a_12420_14488# 0.41329f
C593 a_12754_16434# VDD 0
C594 a_11848_15156# sg13_nor2_1_0.A 0.00241f
C595 adc_start a_16458_14020# 0
C596 sg13_a21oi_1_0.A1 a_15505_16357# 0
C597 timer_done a_13960_4782# 0
C598 a_14246_15234# a_14532_15552# 0.41329f
C599 a_16832_15366# a_16735_15972# 0
C600 a_14820_13735# VDD 0.0085f
C601 a_15217_16349# sg13_o21ai_1_0.B1 0
C602 a_14949_13701# sg13_dfrbpq_1_1.Q 0
C603 a_15051_13844# a_15784_14570# 0
C604 a_12228_13735# sg13_nor2_1_0.B 0
C605 a_14532_15552# sg13_inv_1_1.A 0.01632f
C606 a_15496_16878# sg13_dfrbpq_1_0.CLK 0.00121f
C607 a_13192_12342# sg13_dfrbpq_1_0.CLK 0
C608 a_14248_4688# a_14144_4782# 0.00624f
C609 sg13_nor2b_1_0.Y VDD 0.36901f
C610 a_12134_14922# a_13679_14845# 0
C611 a_12420_14488# a_13297_14837# 0.01835f
C612 a_12394_14452# a_12939_14495# 0.01f
C613 a_12837_14495# a_12708_14909# 0.01562f
C614 sg13_a21oi_1_0.A1 tx_start 0.19049f
C615 a_15872_25498# VDD 0
C616 a_15096_17064# a_14998_16742# 0.00202f
C617 a_14246_15234# a_15791_15311# 0
C618 a_16048_13942# sg13_dfrbpq_1_1.Q 0.00197f
C619 a_13401_14037# a_12459_13844# 0
C620 a_12166_13735# a_11940_14040# 0.0052f
C621 a_12228_13735# a_12357_13701# 0.01562f
C622 a_14340_16000# a_14628_16421# 0.43707f
C623 a_25856_17594# VDD 0.08554f
C624 a_15791_15311# sg13_inv_1_1.A 0.01731f
C625 a_13459_12404# VDD 0.33748f
C626 a_16735_15972# sg13_dfrbpq_1_5.Q 0.04761f
C627 a_12939_14495# a_13936_14726# 0.03061f
C628 a_11464_13644# VDD 0.00177f
C629 a_9920_16426# sg13_dfrbpq_1_0.CLK 0
C630 sg13_and2_1_0.X VDD 0.80231f
C631 a_12166_13735# sg13_inv_1_0.Y 0
C632 a_14532_15552# a_14820_15247# 0.43707f
C633 sg13_inv_1_1.A a_13871_16823# 0
C634 a_14340_16000# sg13_a21oi_1_0.A2 0.00165f
C635 a_13459_12404# a_13105_13799# 0
C636 sg13_buf_1_0.A a_13472_4782# 0.02359f
C637 sg13_buf_1_4.A a_14506_13945# 0
C638 a_14757_16007# sg13_dfrbpq_1_3.Q 0
C639 a_15697_13799# a_15784_14570# 0
C640 sg13_a21oi_1_0.A1 a_14128_16966# 0.0071f
C641 sg13_nor2_1_0.A a_10790_16434# 0.00393f
C642 a_14346_14484# a_14098_14922# 0
C643 a_14998_16742# sg13_dfrbpq_1_6.D 0.10668f
C644 sg13_buf_1_5.X a_14152_10736# 0.28141f
C645 a_17024_13644# sg13_a21o_1_1.A2 0
C646 a_16048_15454# a_15993_15549# 0.00412f
C647 sg13_o21ai_1_0.A1 a_14998_16742# 0.10047f
C648 a_14628_16421# sg13_a21oi_1_0.A2 0
C649 sg13_inv_1_0.Y sg13_dfrbpq_1_1.Q 0.00108f
C650 sg13_o21ai_1_0.B1 a_14314_15964# 0
C651 a_15856_16238# a_15599_16357# 0.34468f
C652 a_13585_14845# sg13_a21oi_1_0.A2 0
C653 sg13_dfrbpq_1_3.D a_14532_15552# 0.04268f
C654 a_14506_15457# a_14949_15213# 0.02242f
C655 a_12652_16119# sg13_dfrbpq_1_4.D 0
C656 sg13_inv_1_0.Y a_13996_14607# 0.01431f
C657 sg13_dfrbpq_1_4.D a_12939_14495# 0
C658 sg13_a21oi_1_0.A1 sg13_dfrbpq_1_0.CLK 0.57077f
C659 sg13_inv_1_1.A a_13777_16823# 0
C660 a_16018_16434# sg13_dfrbpq_1_5.Q 0
C661 sg13_a22oi_1_0.B2 a_14912_16668# 0.00112f
C662 sg13_a21oi_1_0.A1 a_14290_16746# 0
C663 a_11464_13854# VDD 0.15557f
C664 a_12592_16238# sg13_nor2_1_0.Y 0.04449f
C665 a_14152_10736# Timer_en 0.08749f
C666 a_16458_15532# a_16210_15234# 0
C667 a_14757_16007# a_14054_16434# 0.02432f
C668 a_14820_15247# a_14758_15247# 0
C669 a_14949_15213# a_14532_14040# 0
C670 a_15051_15356# sg13_dfrbpq_1_5.Q 0
C671 sg13_dfrbpq_1_3.D a_15791_15311# 0.01921f
C672 a_14532_15552# a_14949_13701# 0
C673 sg13_nor2_1_0.A a_11433_16043# 0
C674 a_15801_16119# sg13_inv_1_0.Y 0.00351f
C675 sg13_dfrbpq_1_0.CLK a_12136_16668# 0.00194f
C676 a_12817_13743# sg13_a21o_1_0.X 0.00118f
C677 sg13_a21oi_1_0.A1 a_11076_16000# 0
C678 a_13029_16725# a_14128_16966# 0
C679 a_13131_16868# a_13871_16823# 0.26905f
C680 sg13_dfrbpq_1_4.D a_13297_14486# 0
C681 a_17696_15366# VDD 0.09234f
C682 uart_en VDD 0.17827f
C683 a_25856_16878# a_25856_17594# 0
C684 a_15993_15549# sg13_dfrbpq_1_0.CLK 0
C685 a_14440_5412# Timer_en 0.00334f
C686 sg13_nor2_1_0.B sg13_nor2_1_0.Y 0.24938f
C687 a_13576_4688# VDD 0.26091f
C688 a_14155_12256# sg13_and2_1_0.X 0.00112f
C689 sg13_a21o_1_0.A2 a_13838_12256# 0
C690 a_14314_15964# a_14346_14484# 0
C691 sg13_dfrbpq_1_3.D a_14758_15247# 0
C692 sg13_nor2_1_0.A a_11654_13722# 0.00114f
C693 adc_en a_14144_4782# 0.00179f
C694 sg13_a21oi_1_0.A1 a_12335_16357# 0
C695 a_14340_16000# VDD 0.10215f
C696 a_13131_16868# a_13489_17042# 0.02138f
C697 a_13029_16725# sg13_dfrbpq_1_0.CLK 0.26754f
C698 sg13_inv_1_1.A a_16108_14037# 0
C699 sg13_inv_1_1.A adc_done 0.00169f
C700 a_14246_15234# sg13_nor2_1_0.B 0
C701 a_13459_12404# a_13480_10830# 0
C702 sg13_a21oi_1_0.A1 a_14188_17061# 0.00134f
C703 a_14506_15457# sg13_dfrbpq_1_0.CLK 0.00419f
C704 a_13960_4572# VDD 0.00206f
C705 a_12838_16759# sg13_dfrbpq_1_0.CLK 0
C706 a_13777_16823# a_13131_16868# 0.00647f
C707 a_25768_14570# VDD 0.15802f
C708 a_14148_16434# sg13_a21oi_1_0.A2 0
C709 a_15697_15311# sg13_dfrbpq_1_5.Q 0
C710 a_13866_14020# a_13679_14845# 0
C711 a_16048_15454# a_15791_13799# 0
C712 a_15791_15311# a_16048_13942# 0
C713 sg13_a21o_1_1.A2 a_16832_15156# 0.00232f
C714 sg13_inv_1_1.A sg13_nor2_1_0.B 0
C715 a_14628_16421# VDD 0.008f
C716 sg13_a22oi_1_0.B2 a_15217_15998# 0
C717 sg13_dfrbpq_1_0.CLK a_10790_16434# 0.0156f
C718 a_13585_14845# VDD 0.00479f
C719 sg13_a22oi_1_0.B2 a_14248_23556# 0
C720 tx_start a_15976_25068# 0
C721 a_12134_14922# a_13996_14607# 0
C722 a_14532_14040# sg13_dfrbpq_1_0.CLK 0.07449f
C723 a_14998_16742# sg13_o21ai_1_0.B1 0.03467f
C724 a_13401_14037# sg13_buf_1_0.A 0
C725 sg13_a21oi_1_0.A2 VDD 2.5718f
C726 a_14532_15552# sg13_inv_1_0.Y 0.4149f
C727 a_14757_16007# sg13_inv_1_1.Y 0
C728 a_16430_14832# a_16051_14746# 0
C729 sg13_dfrbpq_1_3.D a_15051_13844# 0.00277f
C730 a_16294_14484# sg13_a21o_1_1.A2 0.01685f
C731 sg13_dfrbpq_1_0.CLK a_11953_16349# 0.00332f
C732 a_13029_16725# a_12335_16357# 0.00312f
C733 a_12612_17064# a_13002_15996# 0
C734 a_10790_16434# a_11076_16000# 0.41329f
C735 sg13_dfrbpq_1_6.D a_12326_16746# 0.29362f
C736 a_17800_15272# sg13_inv_2_1.A 0.26119f
C737 a_15791_13799# sg13_dfrbpq_1_0.CLK 0.00372f
C738 a_12939_14495# a_13881_14607# 0
C739 a_14054_16434# a_14314_15964# 0.75507f
C740 a_15856_16238# a_15784_14570# 0
C741 a_15791_15311# sg13_inv_1_0.Y 0.13303f
C742 a_14073_17061# sg13_dfrbpq_1_6.D 0
C743 a_14532_14040# a_15409_14018# 0
C744 a_14246_13722# a_14889_14113# 0.00801f
C745 a_14949_13701# a_15051_13844# 0.47622f
C746 a_10790_16434# a_12335_16357# 0
C747 a_11050_15964# a_11595_16007# 0.01f
C748 a_11076_16000# a_11953_16349# 0.01835f
C749 a_11493_16007# a_11364_16421# 0.01562f
C750 sg13_nor2_1_0.A sg13_a21o_1_0.X 0
C751 sg13_inv_1_1.Y a_14098_14922# 0
C752 a_15599_16357# a_16051_14746# 0
C753 reset a_8776_13644# 0.00207f
C754 a_16832_15366# sg13_inv_2_1.A 0.019f
C755 sg13_inv_1_0.Y a_13871_16823# 0.14402f
C756 sg13_dfrbpq_1_3.D sg13_nor2_1_0.B 0
C757 sg13_dfrbpq_1_3.Q sg13_a21o_1_1.A2 0.30602f
C758 a_16832_15366# sg13_a22oi_1_0.B2 0
C759 a_15096_17064# sg13_dfrbpq_1_6.D 0.01075f
C760 a_14758_15247# sg13_inv_1_0.Y 0
C761 a_14148_16434# VDD 0
C762 a_13768_10736# timer_done 0.01199f
C763 sg13_dfrbpq_1_0.CLK a_11654_13722# 0
C764 a_15051_13844# a_16048_13942# 0.02979f
C765 a_14859_16007# a_15801_16119# 0
C766 a_11595_16007# a_12592_16238# 0.03061f
C767 sg13_dfrbpq_1_3.D a_15697_13799# 0
C768 sg13_o21ai_1_0.A1 a_15096_17064# 0.00139f
C769 a_12586_16969# sg13_dfrbpq_1_0.CLK 0
C770 sg13_inv_1_0.Y a_13489_17042# 0.01491f
C771 sg13_inv_2_1.A sg13_dfrbpq_1_5.Q 0.00612f
C772 a_13192_12342# sg13_buf_1_0.A 0.00152f
C773 sg13_nor2b_1_0.Y a_11493_16007# 0.00272f
C774 a_14336_5842# timer_done 0.00106f
C775 a_13777_16823# sg13_inv_1_0.Y 0
C776 sg13_a22oi_1_0.B2 sg13_dfrbpq_1_5.Q 0.3115f
C777 a_13002_15996# a_12754_16434# 0
C778 a_11595_16007# sg13_nor2_1_0.B 0
C779 a_16048_13942# a_16108_14037# 0.01042f
C780 a_15051_13844# a_15409_13743# 0.00104f
C781 a_14949_13701# a_15697_13799# 0.01058f
C782 a_15791_13799# a_16458_14020# 0.0894f
C783 a_14440_5412# a_14248_4688# 0
C784 a_12652_16119# sg13_nor2_1_0.Y 0
C785 a_14757_16007# a_15505_16357# 0.01058f
C786 sg13_nor2_1_0.Y a_12939_14495# 0
C787 sg13_dfrbpq_1_6.D a_12241_16357# 0.00206f
C788 sg13_inv_1_0.Y a_11050_15964# 0.2637f
C789 a_13105_13799# VDD 0.00294f
C790 a_16048_13942# a_15697_13799# 0.008f
C791 a_15051_13844# sg13_inv_1_0.Y 0.42489f
C792 sg13_inv_1_1.Y a_14314_15964# 0.00404f
C793 a_14949_15213# a_14757_16007# 0
C794 sg13_o21ai_1_0.A1 sg13_dfrbpq_1_6.D 0.34452f
C795 sg13_nor2b_1_0.Y a_12136_16878# 0
C796 sg13_nor2_1_0.Y a_13297_14486# 0
C797 a_11848_15366# sg13_nor2b_1_0.Y 0.00444f
C798 sg13_inv_1_0.Y a_12592_16238# 0.12835f
C799 a_12586_16969# a_12335_16357# 0
C800 sg13_a21oi_1_0.A1 a_13499_15996# 0.03306f
C801 sg13_a21oi_1_0.A1 a_13936_14726# 0
C802 uart_busy a_15872_25498# 0.00127f
C803 a_13664_10620# sg13_buf_1_0.A 0.00203f
C804 sg13_nor2_1_0.B a_11940_14040# 0
C805 a_14532_15552# a_14859_16007# 0
C806 a_16108_14037# sg13_inv_1_0.Y 0.01227f
C807 a_14144_23642# tx_start 0
C808 sg13_dfrbpq_1_0.CLK sg13_a21o_1_0.X 0.002f
C809 sg13_a22oi_1_0.B2 a_15872_25498# 0
C810 a_15856_16238# sg13_inv_1_1.A 0.00216f
C811 sg13_inv_1_0.Y sg13_nor2_1_0.B 0.26833f
C812 sg13_a21oi_1_0.A1 a_15599_16357# 0
C813 a_11654_13722# a_12459_13844# 0.097f
C814 a_11940_14040# a_12357_13701# 0.37291f
C815 sg13_buf_1_4.A sg13_inv_1_1.Y 0
C816 sg13_nor2_1_0.B a_13199_13799# 0
C817 a_15688_25154# a_15872_25154# 0.0524f
C818 a_15697_13799# sg13_inv_1_0.Y 0
C819 a_15096_17064# sg13_o21ai_1_0.B1 0
C820 a_13856_25498# VDD 0
C821 a_15784_14570# a_16051_14746# 0.00872f
C822 sg13_inv_1_0.Y a_12357_13701# 0.07392f
C823 a_16735_15972# VDD 0.30448f
C824 a_11654_13722# a_13516_14037# 0
C825 a_11940_14040# a_13456_13942# 0.00242f
C826 a_12357_13701# a_13199_13799# 0.00332f
C827 sg13_a21oi_1_0.A1 sg13_dfrbpq_1_4.D 0.11522f
C828 a_25856_16878# VDD 0.08554f
C829 a_14757_16007# sg13_dfrbpq_1_0.CLK 0.29738f
C830 a_13864_16082# a_12612_17064# 0
C831 a_14155_12256# VDD 0.00172f
C832 sg13_dfrbpq_1_0.CLK a_12708_14909# 0.0025f
C833 a_16458_15532# sg13_dfrbpq_1_3.Q 0.14438f
C834 a_14340_16000# a_14912_16878# 0
C835 wake_up_sg a_10790_16434# 0
C836 sg13_inv_1_0.Y a_13456_13942# 0.1139f
C837 a_14697_16043# a_14054_16434# 0.00801f
C838 clk a_7816_15996# 0.28839f
C839 a_13838_12256# sg13_buf_1_4.A 0.00232f
C840 a_13199_13799# a_13456_13942# 0.34468f
C841 a_15217_16349# sg13_dfrbpq_1_0.CLK 0.00105f
C842 sg13_nor2b_1_0.Y a_11914_13945# 0
C843 a_12592_16238# a_12134_14922# 0
C844 a_13480_10830# VDD 0.13808f
C845 sg13_dfrbpq_1_0.CLK a_14098_14922# 0
C846 sg13_o21ai_1_0.B1 sg13_dfrbpq_1_6.D 0.22379f
C847 a_16210_15234# sg13_dfrbpq_1_3.Q 0
C848 sg13_dfrbpq_1_3.D a_15856_16238# 0
C849 a_14246_13722# a_13679_14845# 0
C850 a_14152_10736# sg13_buf_1_4.A 0.00135f
C851 a_14506_15457# sg13_buf_1_0.A 0
C852 sg13_o21ai_1_0.A1 sg13_o21ai_1_0.B1 0.03551f
C853 a_16018_16434# VDD 0
C854 sg13_inv_1_0.Y a_8776_13644# 0
C855 a_25768_25154# VDD 0.13581f
C856 a_12537_16119# a_12592_16238# 0.00412f
C857 a_12652_16119# a_11595_16007# 0
C858 a_12335_16357# a_12708_14909# 0
C859 a_13029_16725# sg13_dfrbpq_1_4.D 0
C860 sg13_a21o_1_0.X a_12459_13844# 0.00127f
C861 a_14152_5498# VDD 0.1537f
C862 sg13_nor2_1_0.B a_12134_14922# 0.00347f
C863 Timer_en a_13472_4572# 0
C864 sg13_inv_2_1.A a_17696_15366# 0.00301f
C865 wake_up_sg a_11433_16043# 0
C866 a_16266_15996# sg13_dfrbpq_1_5.Q 0.12951f
C867 a_15051_15356# VDD 0.19201f
C868 a_14340_16000# a_14538_17044# 0
C869 a_14532_14040# sg13_buf_1_0.A 0.03105f
C870 sg13_buf_1_5.X sg13_buf_1_0.A 0.00377f
C871 a_15496_16878# a_15680_16878# 0.0524f
C872 sg13_nor2b_1_0.Y a_12420_14488# 0.00199f
C873 sg13_dfrbpq_1_4.D a_10790_16434# 0.28718f
C874 sg13_nor2_1_0.B a_13297_14837# 0
C875 a_14566_16421# sg13_dfrbpq_1_6.D 0
C876 sg13_a22oi_1_0.B2 a_14340_16000# 0.03762f
C877 a_16108_15549# VDD 0.00674f
C878 Timer_en sg13_buf_1_0.A 6.40005f
C879 a_14628_16421# a_14538_17044# 0
C880 sg13_inv_1_0.Y a_12228_14922# 0
C881 sg13_dfrbpq_1_0.CLK a_14314_15964# 0.0201f
C882 sg13_inv_1_1.A a_16051_14746# 0.00355f
C883 sg13_nor2_1_0.B a_12777_14531# 0
C884 sg13_a21oi_1_0.A1 a_13601_16344# 0.01147f
C885 a_12136_16878# sg13_a21oi_1_0.A2 0
C886 sg13_a22oi_1_0.B2 a_14628_16421# 0.00526f
C887 a_14538_17044# sg13_a21oi_1_0.A2 0.00231f
C888 a_15697_15311# VDD 0.0013f
C889 a_12652_16119# sg13_inv_1_0.Y 0.01938f
C890 sg13_inv_1_0.Y a_12939_14495# 0.43355f
C891 a_25672_11546# a_25856_11546# 0.0524f
C892 a_14506_13945# a_14346_14484# 0.00192f
C893 sg13_and2_1_0.X a_13679_14845# 0.00135f
C894 a_9920_16426# a_10024_15996# 0
C895 a_16048_15454# sg13_a21o_1_1.A2 0
C896 sg13_dfrbpq_1_4.D a_11433_16043# 0
C897 a_11654_13722# sg13_buf_1_0.A 0
C898 a_13199_13799# a_12939_14495# 0.00198f
C899 a_14949_15213# a_14998_16742# 0
C900 sg13_a22oi_1_0.B2 sg13_a21oi_1_0.A2 0.00121f
C901 a_15856_16238# sg13_inv_1_0.Y 0.09878f
C902 a_14912_16878# VDD 0.0765f
C903 sg13_inv_1_0.Y a_13297_14486# 0.01788f
C904 a_13768_10736# a_13480_10620# 0
C905 sg13_a21o_1_0.A2 sg13_buf_1_0.A 0.0051f
C906 sg13_buf_1_4.A sg13_dfrbpq_1_0.CLK 0.00113f
C907 a_11493_16007# VDD 0.2548f
C908 sg13_dfrbpq_1_6.D a_14054_16434# 0.00229f
C909 a_16832_15366# sg13_dfrbpq_1_1.Q 0
C910 a_14889_14113# VDD 0
C911 a_14073_17061# sg13_inv_1_1.Y 0
C912 sg13_dfrbpq_1_0.CLK sg13_a21o_1_1.A2 0
C913 sg13_dfrbpq_1_3.D a_16051_14746# 0.17615f
C914 a_12134_14922# a_12228_14922# 0.00716f
C915 adc_start a_16048_13942# 0
C916 a_13002_15996# VDD 0.38576f
C917 sg13_a21oi_1_0.A1 sg13_nor2_1_0.Y 0.03207f
C918 a_12136_16878# VDD 0.15258f
C919 a_14532_14040# a_15784_14570# 0
C920 a_14566_16421# sg13_o21ai_1_0.B1 0
C921 a_17128_13760# VDD 0.23761f
C922 a_14998_16742# sg13_dfrbpq_1_0.CLK 0.00111f
C923 a_14538_17044# VDD 0.38555f
C924 uart_busy VDD 0.1533f
C925 a_13576_4688# a_13960_4782# 0.01f
C926 a_14246_15234# sg13_a21oi_1_0.A1 0
C927 a_12394_14452# a_12708_14909# 0.00463f
C928 a_12420_14488# a_12646_14909# 0.0052f
C929 a_12134_14922# a_12939_14495# 0.097f
C930 a_11848_15366# VDD 0.16361f
C931 a_14144_23986# tx_start 0
C932 a_16735_16388# sg13_inv_1_1.A 0.00132f
C933 sg13_a21o_1_0.X sg13_buf_1_0.A 0.03538f
C934 sg13_inv_2_1.A VDD 0.83109f
C935 a_14437_17878# sg13_a21oi_1_0.A2 0
C936 a_14949_15213# a_15409_15530# 0.01483f
C937 sg13_a21oi_1_0.A1 sg13_inv_1_1.A 0
C938 sg13_nor2b_1_0.Y a_12166_13735# 0
C939 a_15791_13799# a_15784_14570# 0
C940 a_12228_13735# a_11654_13722# 0.31978f
C941 sg13_a22oi_1_0.B2 VDD 2.38189f
C942 sg13_dfrbpq_1_3.Q a_16832_15156# 0.00227f
C943 a_14340_16000# a_13679_14845# 0
C944 a_16840_13644# VDD 0.00177f
C945 a_15801_16119# sg13_dfrbpq_1_5.Q 0
C946 a_12817_14018# VDD 0.00761f
C947 a_12134_14922# a_13297_14486# 0
C948 a_12420_14488# a_13585_14845# 0.43239f
C949 a_13297_14837# a_12939_14495# 0.00104f
C950 a_16048_13942# a_16051_14746# 0.00138f
C951 a_16458_14020# sg13_a21o_1_1.A2 0.00125f
C952 sg13_buf_1_5.X a_13702_12532# 0
C953 a_13401_14037# sg13_inv_1_0.Y 0.00411f
C954 adc_start sg13_inv_1_0.Y 0
C955 sg13_dfrbpq_1_5.Q a_15496_16668# 0.0036f
C956 a_15051_15356# a_16108_15549# 0
C957 sg13_buf_1_0.A a_14248_4688# 0.27925f
C958 a_13029_16725# sg13_nor2_1_0.Y 0.0044f
C959 sg13_dfrbpq_1_6.D sg13_inv_1_1.Y 0
C960 a_12420_14488# sg13_a21oi_1_0.A2 0
C961 a_13866_14020# a_13456_13942# 0.10373f
C962 a_13401_14037# a_13199_13799# 0.00689f
C963 a_14757_16007# a_15599_16357# 0.00307f
C964 a_15993_15549# sg13_inv_1_1.A 0.00183f
C965 a_12838_16759# sg13_nor2_1_0.Y 0
C966 a_13864_16082# a_13585_14845# 0
C967 uart_done a_13856_25154# 0.02302f
C968 a_13679_14845# a_13585_14845# 0.28931f
C969 a_13936_14726# a_14098_14922# 0.00188f
C970 sg13_dfrbpq_1_3.Q a_16294_14484# 0.06804f
C971 a_10790_16434# sg13_nor2_1_0.Y 0
C972 a_15051_15356# a_15697_15311# 0.00647f
C973 sg13_buf_1_0.A a_14144_4572# 0
C974 a_13864_16082# sg13_a21oi_1_0.A2 0.01975f
C975 a_16048_15454# a_16458_15532# 0.10373f
C976 a_17024_13854# sg13_a21o_1_1.A2 0
C977 a_14859_16007# a_15856_16238# 0.03061f
C978 a_14697_16043# sg13_dfrbpq_1_0.CLK 0
C979 sg13_o21ai_1_0.B1 a_14054_16434# 0
C980 a_13679_14845# sg13_a21oi_1_0.A2 0
C981 a_14506_15457# a_14246_15234# 0.75507f
C982 a_14757_16007# sg13_dfrbpq_1_4.D 0
C983 sg13_a21oi_1_0.A1 a_13131_16868# 0.00109f
C984 a_14098_14922# sg13_buf_1_0.A 0
C985 sg13_inv_1_0.Y a_16051_14746# 0.00336f
C986 a_15916_16119# sg13_o21ai_1_0.A1 0
C987 a_14506_15457# sg13_inv_1_1.A 0.01954f
C988 a_15680_16668# sg13_dfrbpq_1_6.D 0
C989 sg13_a21oi_1_0.A1 a_13489_16767# 0
C990 a_11914_13945# VDD 0.09633f
C991 a_15409_15530# sg13_dfrbpq_1_0.CLK 0.00746f
C992 sg13_dfrbpq_1_3.D sg13_a21oi_1_0.A1 0
C993 a_13960_25068# sg13_a21oi_1_0.A2 0.27683f
C994 sg13_inv_2_1.A a_16735_15972# 0.03263f
C995 a_16048_15454# a_16210_15234# 0.00188f
C996 a_14235_17564# sg13_a21oi_1_0.A2 0.19758f
C997 a_14532_15552# sg13_dfrbpq_1_5.Q 0
C998 sg13_o21ai_1_0.A1 a_15680_16668# 0
C999 sg13_a22oi_1_0.B2 a_16735_15972# 0.06687f
C1000 a_12228_13735# sg13_a21o_1_0.X 0.00176f
C1001 sg13_nor2_1_0.A a_12241_16357# 0
C1002 a_14437_17878# VDD 0.00225f
C1003 a_12612_17064# a_13871_16823# 0.01529f
C1004 sg13_nor2_1_0.A sg13_dfrbpq_1_6.D 0
C1005 a_14073_17061# a_14128_16966# 0.00412f
C1006 a_16458_15532# sg13_dfrbpq_1_0.CLK 0.00102f
C1007 a_14152_5842# Timer_en 0.0043f
C1008 a_13192_12342# sg13_inv_1_0.Y 0
C1009 sg13_a21o_1_0.A2 a_13702_12532# 0.01543f
C1010 a_12268_15532# sg13_nor2_1_0.A 0
C1011 a_15791_15311# sg13_dfrbpq_1_5.Q 0.00206f
C1012 sg13_dfrbpq_1_3.D a_15993_15549# 0
C1013 a_14506_15457# a_14820_15247# 0.00463f
C1014 adc_en a_13472_4572# 0
C1015 sg13_a21oi_1_0.A1 a_11595_16007# 0
C1016 Timer_en a_14336_5498# 0.00186f
C1017 a_12420_14488# VDD 0.09197f
C1018 a_16840_13854# VDD 0.12896f
C1019 a_12612_17064# a_13489_17042# 0
C1020 a_12326_16746# sg13_dfrbpq_1_0.CLK 0.00266f
C1021 a_13029_16725# a_13131_16868# 0.47622f
C1022 sg13_inv_1_1.A a_15791_13799# 0
C1023 a_15505_16357# sg13_o21ai_1_0.A1 0.00156f
C1024 a_13960_4782# VDD 0.12486f
C1025 a_13777_16823# a_12612_17064# 0.43239f
C1026 a_13489_16767# a_13029_16725# 0.02396f
C1027 a_25768_14914# VDD 0.0025f
C1028 a_14949_15213# sg13_dfrbpq_1_6.D 0
C1029 a_13866_14020# a_12939_14495# 0
C1030 sg13_nor2_1_0.A a_12297_14113# 0
C1031 a_14949_15213# sg13_o21ai_1_0.A1 0
C1032 a_13864_16082# VDD 0.14373f
C1033 a_12586_16969# sg13_nor2_1_0.Y 0.00153f
C1034 a_13679_14845# VDD 0.20183f
C1035 a_14506_15457# sg13_dfrbpq_1_3.D 0.00465f
C1036 sg13_a22oi_1_0.B2 a_16018_16434# 0
C1037 tx_start a_15688_25498# 0
C1038 a_15051_15356# sg13_inv_2_1.A 0
C1039 adc_en sg13_buf_1_0.A 0.03686f
C1040 a_13960_25068# VDD 0.27901f
C1041 a_15051_15356# sg13_a22oi_1_0.B2 0.00172f
C1042 sg13_dfrbpq_1_4.D a_14314_15964# 0
C1043 a_17800_15272# adc_done 0.25767f
C1044 a_16458_15532# a_16458_14020# 0
C1045 a_14235_17564# VDD 0.29958f
C1046 a_10790_16434# a_10884_16434# 0.00716f
C1047 a_13702_12532# sg13_a21o_1_0.X 0
C1048 sg13_dfrbpq_1_3.D a_14532_14040# 0.00175f
C1049 a_16266_15996# VDD 0.38483f
C1050 sg13_dfrbpq_1_0.CLK a_11302_16421# 0
C1051 a_12612_17064# a_12592_16238# 0
C1052 a_12326_16746# a_12335_16357# 0
C1053 a_16430_14832# sg13_a21o_1_1.A2 0
C1054 sg13_a21oi_1_0.A1 sg13_inv_1_0.Y 0.01437f
C1055 sg13_dfrbpq_1_6.D a_14128_16966# 0.01201f
C1056 sg13_o21ai_1_0.A1 a_14128_16966# 0
C1057 a_14188_17061# a_12326_16746# 0
C1058 a_16108_15549# sg13_a22oi_1_0.B2 0.00104f
C1059 sg13_buf_1_4.A sg13_buf_1_0.A 2.89439f
C1060 a_11848_15156# sg13_inv_1_0.Y 0.0022f
C1061 a_14246_13722# a_15051_13844# 0.097f
C1062 a_14532_14040# a_14949_13701# 0.37291f
C1063 a_12612_17064# sg13_nor2_1_0.B 0
C1064 sg13_dfrbpq_1_0.CLK a_12241_16357# 0.00509f
C1065 a_11050_15964# a_11364_16421# 0.00463f
C1066 a_10790_16434# a_11595_16007# 0.097f
C1067 a_11076_16000# a_11302_16421# 0.0052f
C1068 sg13_dfrbpq_1_3.D a_15791_13799# 0
C1069 sg13_dfrbpq_1_6.D sg13_dfrbpq_1_0.CLK 0.14451f
C1070 sg13_inv_1_0.Y a_12136_16668# 0.00148f
C1071 a_12650_15532# sg13_nor2_1_0.B 0
C1072 a_15697_15311# sg13_inv_2_1.A 0
C1073 a_15993_14037# sg13_dfrbpq_1_0.CLK 0
C1074 a_14290_16746# sg13_dfrbpq_1_6.D 0
C1075 sg13_o21ai_1_0.A1 sg13_dfrbpq_1_0.CLK 0
C1076 a_13864_16426# sg13_a21oi_1_0.A2 0.00434f
C1077 a_15993_15549# sg13_inv_1_0.Y 0.00351f
C1078 a_14246_13722# a_16108_14037# 0
C1079 a_14532_14040# a_16048_13942# 0.00242f
C1080 a_14949_13701# a_15791_13799# 0.00332f
C1081 a_11953_16349# a_11595_16007# 0.00104f
C1082 a_11076_16000# a_12241_16357# 0.43239f
C1083 sg13_dfrbpq_1_3.D a_14758_13735# 0
C1084 a_10790_16434# a_11953_15998# 0
C1085 a_14538_17044# a_14912_16878# 0.01061f
C1086 a_12136_16878# a_11493_16007# 0
C1087 sg13_dfrbpq_1_6.D a_11076_16000# 0.0027f
C1088 sg13_inv_1_0.Y a_13029_16725# 0.03573f
C1089 a_12586_16969# a_13131_16868# 0.01f
C1090 a_13856_25498# a_13960_25068# 0
C1091 a_14506_13945# sg13_dfrbpq_1_0.CLK 0.00212f
C1092 sg13_a22oi_1_0.B2 a_14912_16878# 0.00118f
C1093 a_11848_15366# a_11493_16007# 0.0024f
C1094 a_12838_16759# sg13_inv_1_0.Y 0
C1095 a_14532_14040# a_15409_13743# 0.01835f
C1096 a_15051_13844# a_14820_13735# 0.12701f
C1097 a_15791_13799# a_16048_13942# 0.34468f
C1098 a_12592_16238# a_12754_16434# 0.00188f
C1099 a_12335_16357# a_12241_16357# 0.28931f
C1100 a_14506_15457# sg13_inv_1_0.Y 0.27187f
C1101 a_14949_15213# sg13_o21ai_1_0.B1 0
C1102 sg13_dfrbpq_1_3.Q a_15916_16119# 0
C1103 sg13_dfrbpq_1_6.D a_12335_16357# 0.00371f
C1104 sg13_nor2_1_0.Y a_12708_14909# 0
C1105 sg13_inv_1_0.Y a_10790_16434# 0.11209f
C1106 a_14336_5498# a_14248_4688# 0
C1107 a_12166_13735# VDD 0
C1108 clk VDD 0.65894f
C1109 sg13_buf_1_5.X sg13_inv_1_0.Y 0
C1110 sg13_inv_1_1.Y a_14054_16434# 0.26917f
C1111 a_14532_14040# sg13_inv_1_0.Y 0.38326f
C1112 a_14188_17061# sg13_dfrbpq_1_6.D 0.0018f
C1113 sg13_and2_1_0.X a_15051_13844# 0.00115f
C1114 uart_done tx_start 0.40981f
C1115 a_14757_16007# sg13_inv_1_1.A 0.00313f
C1116 reset a_8968_13760# 0.27187f
C1117 a_12046_15276# a_12268_15532# 0
C1118 sg13_inv_1_0.Y a_11953_16349# 0.00139f
C1119 sg13_inv_2_1.A a_17128_13760# 0
C1120 sg13_nor2b_1_0.Y sg13_nor2_1_0.B 0.19316f
C1121 a_13664_10830# sg13_buf_1_0.A 0.00635f
C1122 a_15791_13799# sg13_inv_1_0.Y 0.13309f
C1123 a_15916_16119# a_14054_16434# 0
C1124 a_13864_16426# VDD 0.0029f
C1125 sg13_a22oi_1_0.B2 uart_busy 0.01152f
C1126 sg13_dfrbpq_1_1.Q VDD 0.78964f
C1127 a_16840_13644# a_17128_13760# 0
C1128 a_16266_15996# a_16018_16434# 0
C1129 sg13_a22oi_1_0.B2 sg13_inv_2_1.A 0.20446f
C1130 sg13_inv_1_1.A a_14098_14922# 0
C1131 sg13_nor2b_1_0.Y a_12357_13701# 0
C1132 sg13_a21oi_1_0.A1 a_14859_16007# 0.00325f
C1133 a_14340_16000# a_13871_16823# 0.00213f
C1134 sg13_inv_1_0.Y a_11433_16043# 0
C1135 a_13996_14607# VDD 0.00816f
C1136 a_11654_13722# a_11940_14040# 0.41329f
C1137 tx_start a_13856_25154# 0
C1138 sg13_o21ai_1_0.B1 sg13_dfrbpq_1_0.CLK 0
C1139 a_14949_15213# sg13_dfrbpq_1_3.Q 0
C1140 a_15976_25068# a_15688_25154# 0.00536f
C1141 sg13_inv_1_0.Y a_11654_13722# 0.1326f
C1142 a_15801_16119# VDD 0
C1143 sg13_and2_1_0.X a_15697_13799# 0
C1144 a_14697_16043# sg13_dfrbpq_1_4.D 0
C1145 a_11654_13722# a_13199_13799# 0
C1146 a_13192_12132# VDD 0.00226f
C1147 a_16048_15454# sg13_dfrbpq_1_3.Q 0.00285f
C1148 a_15496_16668# VDD 0.00217f
C1149 a_12586_16969# sg13_inv_1_0.Y 0.2481f
C1150 sg13_dfrbpq_1_0.CLK a_12837_14495# 0.28366f
C1151 sg13_a21o_1_0.A2 sg13_inv_1_0.Y 0
C1152 sg13_dfrbpq_1_3.D a_14757_16007# 0
C1153 sg13_dfrbpq_1_0.CLK a_16294_14484# 0
C1154 sg13_buf_1_5.X timer_done 0.04183f
C1155 sg13_inv_1_0.Y a_11748_13722# 0
C1156 a_13871_16823# sg13_a21oi_1_0.A2 0.01596f
C1157 a_13702_12532# sg13_buf_1_4.A 0.08185f
C1158 a_13459_12404# a_13456_13942# 0
C1159 a_13768_10736# VDD 0.24991f
C1160 a_9920_16082# VDD 0.09231f
C1161 a_14246_15234# a_14314_15964# 0
C1162 sg13_dfrbpq_1_0.CLK a_14346_14484# 0.00188f
C1163 sg13_inv_1_1.A a_14314_15964# 0.00181f
C1164 a_16735_15972# sg13_dfrbpq_1_1.Q 0
C1165 a_13489_17042# sg13_a21oi_1_0.A2 0.00419f
C1166 timer_done Timer_en 2.27389f
C1167 adc_done a_17696_15366# 0.02303f
C1168 sg13_dfrbpq_1_3.Q sg13_dfrbpq_1_0.CLK 0.02791f
C1169 a_12335_16357# a_12837_14495# 0.00109f
C1170 sg13_a21o_1_0.X a_11940_14040# 0.00907f
C1171 a_14336_5842# VDD 0.00255f
C1172 a_13777_16823# sg13_a21oi_1_0.A2 0.0141f
C1173 a_15856_16238# sg13_dfrbpq_1_5.Q 0.0065f
C1174 a_14532_15552# VDD 0.09587f
C1175 a_16840_13854# a_17128_13760# 0.00536f
C1176 a_14128_16966# a_14054_16434# 0
C1177 sg13_nor2b_1_0.Y a_12228_14922# 0
C1178 sg13_inv_1_0.Y sg13_a21o_1_0.X 0.15319f
C1179 adc_done a_25768_14570# 0.00255f
C1180 sg13_a21o_1_0.X a_13199_13799# 0
C1181 a_15791_15311# VDD 0.17635f
C1182 sg13_inv_1_1.A sg13_buf_1_4.A 0
C1183 clk_gating_en sg13_buf_1_0.A 0.0021f
C1184 a_13618_13722# sg13_buf_1_0.A 0
C1185 sg13_dfrbpq_1_0.CLK a_14054_16434# 0.02387f
C1186 a_17800_15272# adc_start 0
C1187 a_12459_13844# a_12837_14495# 0
C1188 a_13871_16823# VDD 0.18863f
C1189 sg13_a22oi_1_0.B2 a_13864_16082# 0
C1190 a_14757_16007# sg13_inv_1_0.Y 0.0418f
C1191 sg13_inv_1_1.A sg13_a21o_1_1.A2 0.01042f
C1192 a_14758_15247# VDD 0
C1193 sg13_dfrbpq_1_3.Q a_16458_14020# 0
C1194 sg13_dfrbpq_1_3.D a_14314_15964# 0.00107f
C1195 a_14235_17564# a_14538_17044# 0
C1196 a_15599_16357# sg13_o21ai_1_0.A1 0.00137f
C1197 sg13_inv_1_0.Y a_12708_14909# 0.01117f
C1198 sg13_dfrbpq_1_4.D a_12241_16357# 0
C1199 sg13_inv_1_0.Y a_8968_13760# 0
C1200 a_13489_17042# VDD 0.00737f
C1201 sg13_a22oi_1_0.B2 a_14235_17564# 0
C1202 sg13_a22oi_1_0.B2 a_16266_15996# 0.01551f
C1203 sg13_dfrbpq_1_6.D sg13_dfrbpq_1_4.D 0
C1204 a_13777_16823# VDD 0.00374f
C1205 sg13_inv_1_0.Y a_14098_14922# 0
C1206 a_13768_10736# a_13480_10830# 0.00536f
C1207 sg13_a21oi_1_0.A1 a_14912_16668# 0.00305f
C1208 a_14144_17594# sg13_o21ai_1_0.B1 0
C1209 a_12817_13743# sg13_dfrbpq_1_0.CLK 0.00155f
C1210 a_12268_15532# sg13_dfrbpq_1_4.D 0
C1211 a_14506_13945# sg13_buf_1_0.A 0.03218f
C1212 a_14128_16966# sg13_inv_1_1.Y 0
C1213 a_11050_15964# VDD 0.10011f
C1214 a_8968_13760# a_8776_13854# 0.01209f
C1215 a_15051_13844# VDD 0.19677f
C1216 a_16210_13722# a_16458_14020# 0
C1217 a_12592_16238# VDD 0.16101f
C1218 sg13_dfrbpq_1_0.CLK sg13_inv_1_1.Y 0.08915f
C1219 sg13_dfrbpq_1_3.D sg13_a21o_1_1.A2 0.00223f
C1220 timer_done a_14248_4688# 0.04818f
C1221 a_16108_14037# VDD 0.00683f
C1222 adc_done VDD 1.70252f
C1223 a_14949_15213# a_15505_16357# 0
C1224 a_14248_4688# a_14632_4688# 0.0015f
C1225 a_13576_4688# a_13472_4782# 0.00624f
C1226 a_12134_14922# a_12708_14909# 0.31978f
C1227 a_12394_14452# a_12837_14495# 0.02242f
C1228 sg13_nor2_1_0.B VDD 0.61243f
C1229 a_14697_16043# sg13_inv_1_1.A 0
C1230 a_15916_16119# sg13_dfrbpq_1_0.CLK 0.00214f
C1231 a_14246_15234# a_15409_15530# 0
C1232 a_14532_15552# a_15051_15356# 0.34114f
C1233 sg13_inv_1_0.Y a_14314_15964# 0.26514f
C1234 timer_done a_14144_4572# 0.00139f
C1235 a_15697_13799# VDD 0.00289f
C1236 a_14248_23556# sg13_a21oi_1_0.A1 0.28481f
C1237 a_14235_17564# a_14437_17878# 0.01117f
C1238 a_13499_15996# a_12837_14495# 0
C1239 a_16430_14832# a_16294_14484# 0
C1240 a_15409_15530# sg13_inv_1_1.A 0.00263f
C1241 a_12420_14488# a_13679_14845# 0.01529f
C1242 a_12837_14495# a_13936_14726# 0
C1243 a_12708_14909# a_13297_14837# 0
C1244 a_12357_13701# VDD 0.25525f
C1245 a_15872_25154# VDD 0.06317f
C1246 sg13_buf_1_5.X a_14061_12256# 0.26753f
C1247 sg13_dfrbpq_1_5.Q a_15496_16878# 0.00376f
C1248 sg13_dfrbpq_1_6.D a_13601_16344# 0
C1249 a_12326_16746# sg13_nor2_1_0.Y 0.0022f
C1250 a_14949_15213# a_16048_15454# 0
C1251 a_15051_15356# a_15791_15311# 0.26905f
C1252 a_14340_16000# a_15856_16238# 0.00139f
C1253 a_14757_16007# a_14859_16007# 0.47795f
C1254 a_17128_13760# sg13_dfrbpq_1_1.Q 0.28934f
C1255 a_12817_13743# a_12459_13844# 0.00104f
C1256 a_13105_13799# a_12357_13701# 0.01058f
C1257 a_13864_16082# a_13679_14845# 0
C1258 a_16458_15532# sg13_inv_1_1.A 0.01694f
C1259 a_8968_13760# sg13_buf_1_6.X 0.24652f
C1260 sg13_nor2_1_0.A sg13_dfrbpq_1_0.CLK 0.04368f
C1261 a_12837_14495# sg13_buf_1_0.A 0
C1262 a_13936_14726# a_14346_14484# 0.10373f
C1263 a_12939_14495# a_13585_14845# 0.00647f
C1264 a_13456_13942# VDD 0.16565f
C1265 sg13_dfrbpq_1_3.Q a_16430_14832# 0.002f
C1266 sg13_inv_2_1.A sg13_dfrbpq_1_1.Q 0.01069f
C1267 sg13_buf_1_4.A sg13_inv_1_0.Y 0.02045f
C1268 a_15791_15311# a_16108_15549# 0.00247f
C1269 sg13_buf_1_0.A a_14144_4782# 0.02493f
C1270 a_14532_15552# a_15697_15311# 0.43239f
C1271 a_14949_15213# a_15409_15255# 0.02396f
C1272 sg13_a22oi_1_0.B2 sg13_dfrbpq_1_1.Q 0
C1273 sg13_buf_1_4.A a_13199_13799# 0.00147f
C1274 a_13105_13799# a_13456_13942# 0.008f
C1275 a_15217_16349# a_14859_16007# 0.00104f
C1276 a_12939_14495# sg13_a21oi_1_0.A2 0
C1277 a_15505_16357# sg13_dfrbpq_1_0.CLK 0.0023f
C1278 sg13_a21oi_1_0.A1 a_12612_17064# 0.00519f
C1279 a_16210_15234# sg13_inv_1_1.A 0
C1280 sg13_nor2_1_0.A a_11076_16000# 0.00133f
C1281 a_16840_13644# sg13_dfrbpq_1_1.Q 0.00624f
C1282 sg13_dfrbpq_1_4.D a_12837_14495# 0
C1283 a_14346_14484# sg13_buf_1_0.A 0.11665f
C1284 a_15680_16878# sg13_dfrbpq_1_6.D 0.00205f
C1285 sg13_inv_1_0.Y sg13_a21o_1_1.A2 0
C1286 a_14949_15213# sg13_dfrbpq_1_0.CLK 0.28261f
C1287 a_8776_13644# VDD 0.00177f
C1288 adc_done a_25856_16878# 0
C1289 a_15791_15311# a_15697_15311# 0.28931f
C1290 a_15599_16357# sg13_dfrbpq_1_3.Q 0.00253f
C1291 sg13_o21ai_1_0.A1 a_15680_16878# 0.00348f
C1292 sg13_a22oi_1_0.B2 a_15801_16119# 0
C1293 sg13_dfrbpq_1_3.D a_15409_15530# 0
C1294 a_14506_15457# a_14889_15625# 0.00333f
C1295 a_12326_16746# a_12420_16746# 0.00716f
C1296 sg13_nor2_1_0.A a_12335_16357# 0
C1297 a_16735_16388# sg13_dfrbpq_1_5.Q 0.00467f
C1298 a_16048_15454# sg13_dfrbpq_1_0.CLK 0.00164f
C1299 sg13_a22oi_1_0.B2 a_15496_16668# 0.00389f
C1300 a_14998_16742# sg13_inv_1_0.Y 0
C1301 sg13_a21oi_1_0.A1 sg13_dfrbpq_1_5.Q 0
C1302 sg13_a21o_1_0.A2 a_14061_12256# 0.00359f
C1303 a_13459_12404# a_13192_12342# 0.00872f
C1304 timer_done adc_en 0
C1305 a_15051_15356# a_15051_13844# 0
C1306 a_12046_15276# sg13_nor2_1_0.A 0.27095f
C1307 a_13499_15996# a_14054_16434# 0.00243f
C1308 sg13_dfrbpq_1_6.D sg13_nor2_1_0.Y 0.00217f
C1309 sg13_dfrbpq_1_3.D a_16458_15532# 0.00156f
C1310 sg13_dfrbpq_1_0.CLK a_14128_16966# 0
C1311 a_12228_14922# VDD 0
C1312 a_12612_17064# a_13029_16725# 0.37291f
C1313 a_12326_16746# a_13131_16868# 0.097f
C1314 a_15409_15255# sg13_dfrbpq_1_0.CLK 0.00635f
C1315 a_12268_15532# sg13_nor2_1_0.Y 0
C1316 a_14290_16746# a_14128_16966# 0.00188f
C1317 a_14073_17061# a_13131_16868# 0
C1318 a_12838_16759# a_12612_17064# 0.0052f
C1319 a_12900_16759# a_13029_16725# 0.01562f
C1320 a_13472_4782# VDD 0.07977f
C1321 a_15599_16357# a_14054_16434# 0
C1322 a_14859_16007# a_14314_15964# 0.01f
C1323 sg13_nor2_1_0.A a_12459_13844# 0
C1324 timer_done sg13_buf_1_4.A 0.00488f
C1325 sg13_a21oi_1_0.A1 a_12754_16434# 0
C1326 a_14246_15234# sg13_o21ai_1_0.A1 0
C1327 a_12652_16119# VDD 0.00648f
C1328 sg13_dfrbpq_1_3.D a_16210_15234# 0
C1329 a_12900_16759# a_12838_16759# 0
C1330 sg13_inv_1_1.A sg13_dfrbpq_1_6.D 0
C1331 adc_start a_25768_14570# 0.00173f
C1332 sg13_inv_1_1.A a_15993_14037# 0
C1333 a_12939_14495# VDD 0.20221f
C1334 sg13_inv_1_1.A sg13_o21ai_1_0.A1 0
C1335 a_14532_15552# sg13_inv_2_1.A 0
C1336 a_25768_4572# VDD 0.00121f
C1337 a_14532_15552# sg13_a22oi_1_0.B2 0
C1338 sg13_dfrbpq_1_4.D a_14054_16434# 0.00212f
C1339 a_15697_15311# a_15051_13844# 0
C1340 a_15856_16238# VDD 0.16243f
C1341 a_25768_23642# VDD 0.15447f
C1342 a_14061_12256# sg13_a21o_1_0.X 0
C1343 a_13297_14486# VDD 0.00826f
C1344 sg13_dfrbpq_1_0.CLK a_11076_16000# 0.10773f
C1345 a_12326_16746# a_11595_16007# 0
C1346 sg13_nor2b_1_0.Y a_11848_15156# 0.00418f
C1347 a_14697_16043# sg13_inv_1_0.Y 0
C1348 sg13_dfrbpq_1_6.D a_12420_16746# 0
C1349 a_16840_13854# sg13_dfrbpq_1_1.Q 0.03283f
C1350 a_15791_15311# sg13_inv_2_1.A 0.00212f
C1351 a_14188_17061# a_14128_16966# 0.01042f
C1352 a_14538_17044# a_13871_16823# 0.0894f
C1353 a_15409_14018# sg13_dfrbpq_1_0.CLK 0.00525f
C1354 a_15791_15311# sg13_a22oi_1_0.B2 0.00161f
C1355 a_12817_13743# sg13_buf_1_0.A 0
C1356 a_15409_15530# sg13_inv_1_0.Y 0.01621f
C1357 sg13_nor2b_1_0.Y a_12136_16668# 0
C1358 a_15680_16878# sg13_o21ai_1_0.B1 0
C1359 a_14820_15247# sg13_o21ai_1_0.A1 0
C1360 a_10790_16434# a_11364_16421# 0.31978f
C1361 a_11050_15964# a_11493_16007# 0.02242f
C1362 a_13499_15996# sg13_inv_1_1.Y 0.00659f
C1363 a_14246_13722# a_14532_14040# 0.41329f
C1364 sg13_dfrbpq_1_0.CLK a_12335_16357# 0.01736f
C1365 sg13_inv_1_1.Y a_13936_14726# 0
C1366 a_13679_14845# a_13996_14607# 0.00247f
C1367 a_12586_16969# a_12969_17137# 0.00333f
C1368 sg13_dfrbpq_1_6.D a_13131_16868# 0.02198f
C1369 a_14340_16000# a_15496_16878# 0
C1370 a_16458_14020# sg13_dfrbpq_1_0.CLK 0
C1371 sg13_o21ai_1_0.A1 a_13131_16868# 0
C1372 a_13489_16767# sg13_dfrbpq_1_6.D 0.00259f
C1373 a_16458_15532# sg13_inv_1_0.Y 0
C1374 a_16266_15996# sg13_dfrbpq_1_1.Q 0
C1375 sg13_dfrbpq_1_3.Q a_15784_14570# 0
C1376 a_12046_15276# sg13_dfrbpq_1_0.CLK 0
C1377 a_14246_13722# a_15791_13799# 0
C1378 a_11493_16007# a_12592_16238# 0
C1379 a_11364_16421# a_11953_16349# 0
C1380 a_11076_16000# a_12335_16357# 0.01529f
C1381 sg13_dfrbpq_1_3.D a_15993_14037# 0
C1382 sg13_inv_1_1.Y sg13_buf_1_0.A 0
C1383 sg13_dfrbpq_1_3.D sg13_o21ai_1_0.A1 0
C1384 sg13_inv_1_0.Y a_12326_16746# 0.08895f
C1385 a_12586_16969# a_12612_17064# 0.36952f
C1386 a_12046_15276# a_11076_16000# 0
C1387 sg13_nor2_1_0.A a_12394_14452# 0
C1388 a_17024_13854# sg13_dfrbpq_1_0.CLK 0
C1389 sg13_dfrbpq_1_0.CLK a_12459_13844# 0.03872f
C1390 a_12900_16759# a_12586_16969# 0.00463f
C1391 a_14073_17061# sg13_inv_1_0.Y 0.00351f
C1392 a_14532_14040# a_14820_13735# 0.43707f
C1393 wake_up_sg sg13_nor2_1_0.A 0.0276f
C1394 a_11493_16007# sg13_nor2_1_0.B 0.0019f
C1395 sg13_dfrbpq_1_4.D sg13_inv_1_1.Y 0
C1396 a_15599_16357# a_15916_16119# 0.00247f
C1397 a_12592_16238# a_13002_15996# 0.10373f
C1398 a_11595_16007# a_12241_16357# 0.00647f
C1399 sg13_dfrbpq_1_3.Q a_17006_16388# 0.00818f
C1400 sg13_dfrbpq_1_3.D a_14506_13945# 0.00131f
C1401 sc_en a_14248_4688# 0
C1402 sg13_nor2_1_0.Y a_12837_14495# 0
C1403 sg13_dfrbpq_1_6.D a_11595_16007# 0
C1404 sg13_inv_1_1.A sg13_o21ai_1_0.B1 0
C1405 sg13_inv_1_1.A a_16832_15156# 0
C1406 a_13401_14037# VDD 0
C1407 adc_start VDD 1.54847f
C1408 a_13838_12256# sg13_buf_1_0.A 0
C1409 sg13_dfrbpq_1_0.CLK a_13516_14037# 0.00414f
C1410 a_13002_15996# sg13_nor2_1_0.B 0.11615f
C1411 a_16048_13942# a_15993_14037# 0.00412f
C1412 sg13_buf_1_5.X sg13_and2_1_0.X 0.01806f
C1413 sg13_and2_1_0.X a_14532_14040# 0.05365f
C1414 a_14506_13945# a_14949_13701# 0.02242f
C1415 a_14757_16007# a_15217_15998# 0.01483f
C1416 sg13_inv_1_0.Y a_11302_16421# 0
C1417 a_12228_13735# a_12817_13743# 0
C1418 a_13866_14020# sg13_buf_1_4.A 0.12094f
C1419 sg13_a21oi_1_0.A1 a_14340_16000# 0.0382f
C1420 a_14144_17594# a_14128_16966# 0
C1421 sg13_inv_2_1.A adc_done 0.23942f
C1422 a_14152_10736# sg13_buf_1_0.A 0
C1423 a_14820_13735# a_14758_13735# 0
C1424 a_13618_13722# sg13_inv_1_0.Y 0
C1425 sg13_inv_1_1.A a_16294_14484# 0.00138f
C1426 sg13_and2_1_0.X a_15791_13799# 0
C1427 a_17800_15272# a_17696_15156# 0
C1428 a_13618_13722# a_13199_13799# 0.00174f
C1429 a_15856_16238# a_16018_16434# 0.00188f
C1430 a_15599_16357# a_15505_16357# 0.28931f
C1431 a_16051_14746# VDD 0.33625f
C1432 sg13_inv_1_0.Y a_12241_16357# 0.00979f
C1433 sg13_a21oi_1_0.A1 a_14628_16421# 0.01928f
C1434 a_14248_23556# a_14144_23642# 0.00624f
C1435 a_25768_25154# a_25768_23642# 0
C1436 sg13_nor2b_1_0.Y a_11654_13722# 0
C1437 uart_busy a_15872_25154# 0.02302f
C1438 sg13_nor2_1_0.B a_12817_14018# 0
C1439 sg13_nor2_1_0.A sg13_dfrbpq_1_4.D 0.11629f
C1440 a_14440_5412# sg13_buf_1_0.A 0.25844f
C1441 sg13_inv_1_0.Y sg13_dfrbpq_1_6.D 0.13773f
C1442 sg13_a21oi_1_0.A1 a_13585_14845# 0
C1443 a_15872_25498# a_15976_25068# 0
C1444 a_14949_15213# a_15599_16357# 0
C1445 a_15051_15356# a_15856_16238# 0
C1446 a_15993_14037# sg13_inv_1_0.Y 0.00351f
C1447 a_12268_15532# sg13_inv_1_0.Y 0
C1448 sg13_dfrbpq_1_3.D sg13_o21ai_1_0.B1 0
C1449 sg13_o21ai_1_0.A1 sg13_inv_1_0.Y 0
C1450 sg13_and2_1_0.X a_14758_13735# 0
C1451 sg13_dfrbpq_1_3.D a_16832_15156# 0
C1452 sg13_a22oi_1_0.B2 a_15872_25154# 0
C1453 sg13_dfrbpq_1_3.Q sg13_inv_1_1.A 0.48813f
C1454 sg13_a21oi_1_0.A1 sg13_a21oi_1_0.A2 0.93858f
C1455 a_13864_16082# a_13871_16823# 0
C1456 a_12357_13701# a_12817_14018# 0.01483f
C1457 a_11654_13722# a_11464_13644# 0.00404f
C1458 a_13192_12342# VDD 0.16299f
C1459 a_15496_16878# VDD 0.12716f
C1460 sg13_dfrbpq_1_0.CLK a_12394_14452# 0.00219f
C1461 a_16048_15454# a_15599_16357# 0.00123f
C1462 a_15791_15311# a_16266_15996# 0.00159f
C1463 wake_up_sg sg13_dfrbpq_1_0.CLK 0.34463f
C1464 a_13601_16344# sg13_inv_1_1.Y 0
C1465 a_14506_13945# sg13_inv_1_0.Y 0.26528f
C1466 a_13459_12404# sg13_a21o_1_0.A2 0.00148f
C1467 sg13_inv_1_0.Y a_12297_14113# 0.00108f
C1468 a_14061_12256# sg13_buf_1_4.A 0.16354f
C1469 a_12459_13844# a_13516_14037# 0
C1470 a_13499_15996# sg13_dfrbpq_1_0.CLK 0.0344f
C1471 a_14235_17564# a_13871_16823# 0.00163f
C1472 sg13_dfrbpq_1_0.CLK a_13936_14726# 0.00361f
C1473 a_9920_16426# VDD 0
C1474 a_25672_11546# VDD 0.13452f
C1475 a_13864_16082# a_13777_16823# 0
C1476 wake_up_sg a_11076_16000# 0
C1477 a_14757_16007# sg13_dfrbpq_1_5.Q 0
C1478 a_15697_15311# a_15856_16238# 0
C1479 sg13_nor2_1_0.B a_11914_13945# 0
C1480 sg13_dfrbpq_1_3.D a_14346_14484# 0.00532f
C1481 sg13_inv_1_1.A a_14054_16434# 0.00301f
C1482 Timer_en uart_en 0.00128f
C1483 a_12228_13735# sg13_nor2_1_0.A 0
C1484 sg13_a21oi_1_0.A1 a_14148_16434# 0
C1485 a_13029_16725# sg13_a21oi_1_0.A2 0.03181f
C1486 Timer_en a_13576_4688# 0.00441f
C1487 clk_gating_en a_14632_4688# 0.24489f
C1488 a_15599_16357# sg13_dfrbpq_1_0.CLK 0.0066f
C1489 a_13664_10620# VDD 0
C1490 a_12592_16238# a_12420_14488# 0
C1491 a_12335_16357# a_12394_14452# 0
C1492 a_11464_13854# a_11654_13722# 0.00201f
C1493 a_11914_13945# a_12357_13701# 0.02242f
C1494 sg13_dfrbpq_1_0.CLK sg13_buf_1_0.A 0.0292f
C1495 a_15217_16349# sg13_dfrbpq_1_5.Q 0
C1496 sg13_dfrbpq_1_3.D sg13_dfrbpq_1_3.Q 0.05039f
C1497 a_16735_16388# VDD 0
C1498 a_14998_16742# a_14912_16668# 0.00206f
C1499 sg13_inv_1_0.Y a_9728_13644# 0
C1500 a_13459_12404# sg13_a21o_1_0.X 0.18127f
C1501 sg13_nor2_1_0.B a_12420_14488# 0.00895f
C1502 Timer_en a_13960_4572# 0.00685f
C1503 sg13_a21oi_1_0.A1 VDD 2.24173f
C1504 sg13_dfrbpq_1_0.CLK sg13_dfrbpq_1_4.D 0.91997f
C1505 sg13_a21o_1_0.X a_11464_13644# 0.00444f
C1506 sg13_and2_1_0.X sg13_a21o_1_0.X 0
C1507 adc_done a_25768_14914# 0.00188f
C1508 a_11848_15156# VDD 0.00181f
C1509 sg13_o21ai_1_0.B1 sg13_inv_1_0.Y 0.00118f
C1510 a_15505_16357# a_15784_14570# 0
C1511 a_13702_12532# a_13838_12256# 0
C1512 sg13_dfrbpq_1_4.D a_11076_16000# 0.0185f
C1513 a_11940_14040# a_12837_14495# 0
C1514 a_13131_16868# a_14054_16434# 0
C1515 a_12136_16668# VDD 0.00121f
C1516 a_14859_16007# sg13_dfrbpq_1_6.D 0.00263f
C1517 a_14949_15213# a_15784_14570# 0.00104f
C1518 a_14246_15234# sg13_inv_1_1.Y 0.02997f
C1519 sg13_dfrbpq_1_3.D a_14054_16434# 0
C1520 a_15993_15549# VDD 0
C1521 a_14859_16007# sg13_o21ai_1_0.A1 0
C1522 sg13_inv_1_0.Y a_12837_14495# 0.04713f
C1523 sg13_inv_1_1.A sg13_inv_1_1.Y 0.11473f
C1524 a_13456_13942# a_12420_14488# 0
C1525 a_13199_13799# a_12837_14495# 0.00173f
C1526 sg13_dfrbpq_1_4.D a_12335_16357# 0.00886f
C1527 a_13029_16725# VDD 0.23908f
C1528 sg13_a22oi_1_0.B2 a_15856_16238# 0.01305f
C1529 a_15791_15311# sg13_dfrbpq_1_1.Q 0.00254f
C1530 a_14566_16421# sg13_inv_1_0.Y 0
C1531 a_11464_13854# sg13_a21o_1_0.X 0.03327f
C1532 a_14340_15234# sg13_inv_1_1.Y 0
C1533 a_15505_16357# a_15680_16878# 0
C1534 sg13_inv_1_0.Y a_14346_14484# 0.01923f
C1535 a_14506_15457# VDD 0.09995f
C1536 a_12838_16759# VDD 0
C1537 a_12228_13735# sg13_dfrbpq_1_0.CLK 0
C1538 a_12046_15276# sg13_dfrbpq_1_4.D 0.00173f
C1539 a_10024_15996# sg13_nor2_1_0.A 0.24593f
C1540 a_17800_15272# sg13_a21o_1_1.A2 0.00112f
C1541 a_12459_13844# sg13_buf_1_0.A 0
C1542 sg13_inv_1_1.A a_15916_16119# 0.00137f
C1543 a_16735_16388# a_16735_15972# 0
C1544 a_10790_16434# VDD 0.78695f
C1545 a_12586_16969# sg13_a21oi_1_0.A2 0.00171f
C1546 sg13_dfrbpq_1_3.Q sg13_inv_1_0.Y 0.00177f
C1547 sg13_nor2_1_0.A sg13_nor2_1_0.Y 0.0898f
C1548 sg13_buf_1_5.X VDD 0.94285f
C1549 a_14532_14040# VDD 0.09642f
C1550 a_15697_15311# a_16051_14746# 0
C1551 a_16832_15366# sg13_a21o_1_1.A2 0.00285f
C1552 a_13516_14037# sg13_buf_1_0.A 0
C1553 sg13_dfrbpq_1_0.CLK a_15784_14570# 0.00697f
C1554 a_11953_16349# VDD 0
C1555 a_16210_13722# a_16048_13942# 0.00188f
C1556 a_13866_14020# a_13618_13722# 0
C1557 sg13_buf_1_4.A a_14246_13722# 0.03688f
C1558 sg13_dfrbpq_1_0.CLK a_13601_16344# 0.00152f
C1559 a_13131_16868# sg13_inv_1_1.Y 0
C1560 sg13_inv_1_1.A sg13_nor2_1_0.A 0.00111f
C1561 uart_en a_14248_4688# 0.24499f
C1562 sg13_dfrbpq_1_0.CLK a_13881_14607# 0.00108f
C1563 a_15791_13799# VDD 0.18497f
C1564 sg13_buf_1_6.X a_9728_13644# 0.00121f
C1565 a_14152_5842# a_14440_5412# 0
C1566 Timer_en VDD 0.94498f
C1567 sg13_dfrbpq_1_3.D sg13_inv_1_1.Y 0.05216f
C1568 a_13576_4688# a_14248_4688# 0
C1569 a_12134_14922# a_12837_14495# 0.02432f
C1570 adc_start a_17128_13760# 0.24584f
C1571 a_11433_16043# VDD 0
C1572 sg13_dfrbpq_1_5.Q sg13_a21o_1_1.A2 0.00349f
C1573 sg13_buf_1_4.A a_14340_13722# 0
C1574 sg13_inv_1_0.Y a_14054_16434# 0.12637f
C1575 a_14440_5412# a_14336_5498# 0.00617f
C1576 a_14246_15234# a_14949_15213# 0.02454f
C1577 timer_done a_14144_4782# 0.00116f
C1578 sg13_a21oi_1_0.A1 a_16018_16434# 0
C1579 a_14758_13735# VDD 0
C1580 a_14144_23986# a_14248_23556# 0
C1581 a_14859_16007# sg13_o21ai_1_0.B1 0
C1582 a_14340_16000# a_14757_16007# 0.37384f
C1583 a_15051_13844# sg13_dfrbpq_1_1.Q 0
C1584 a_14248_4688# a_13960_4572# 0
C1585 a_14949_15213# sg13_inv_1_1.A 0.01628f
C1586 sg13_inv_2_1.A adc_start 0
C1587 a_12646_14909# a_12708_14909# 0
C1588 a_12837_14495# a_13297_14837# 0.02396f
C1589 a_12420_14488# a_12939_14495# 0.34102f
C1590 a_11654_13722# VDD 0.78247f
C1591 a_15976_25068# VDD 0.24955f
C1592 sg13_dfrbpq_1_5.Q a_14998_16742# 0
C1593 a_14532_15552# a_15791_15311# 0.01529f
C1594 a_16840_13644# adc_start 0.00192f
C1595 a_16108_14037# sg13_dfrbpq_1_1.Q 0
C1596 a_12817_13743# a_11940_14040# 0.01835f
C1597 a_12228_13735# a_12459_13844# 0.12701f
C1598 a_13866_14020# a_14506_13945# 0
C1599 a_14340_16000# a_15217_16349# 0.01835f
C1600 a_14757_16007# a_14628_16421# 0.01562f
C1601 a_12586_16969# VDD 0.09717f
C1602 sg13_a21o_1_0.A2 VDD 0.44683f
C1603 a_16048_15454# sg13_inv_1_1.A 0.0143f
C1604 a_13864_16082# a_12939_14495# 0
C1605 a_11748_13722# VDD 0
C1606 a_10024_15996# sg13_dfrbpq_1_0.CLK 0.01283f
C1607 a_12420_14488# a_13297_14486# 0
C1608 a_12939_14495# a_13679_14845# 0.26905f
C1609 sg13_buf_1_5.X a_14155_12256# 0.01071f
C1610 a_12817_13743# sg13_inv_1_0.Y 0.00227f
C1611 a_14532_15552# a_14758_15247# 0.0052f
C1612 sg13_inv_1_1.A a_14128_16966# 0
C1613 a_15051_15356# a_15993_15549# 0
C1614 a_14949_15213# a_14820_15247# 0.01562f
C1615 a_14757_16007# sg13_a21oi_1_0.A2 0
C1616 a_13459_12404# sg13_buf_1_4.A 0.01282f
C1617 sg13_buf_1_4.A sg13_and2_1_0.X 0.15615f
C1618 sg13_dfrbpq_1_0.CLK sg13_nor2_1_0.Y 0.14088f
C1619 a_14628_16421# a_15217_16349# 0
C1620 sg13_a22oi_1_0.B2 a_16051_14746# 0
C1621 a_15409_15255# sg13_inv_1_1.A 0
C1622 a_13585_14845# a_14098_14922# 0
C1623 a_13936_14726# sg13_buf_1_0.A 0.00128f
C1624 wake_up_sg sg13_dfrbpq_1_4.D 0.00922f
C1625 a_14246_15234# sg13_dfrbpq_1_0.CLK 0.00826f
C1626 a_14912_16668# sg13_dfrbpq_1_6.D 0
C1627 a_14144_23642# sg13_a21oi_1_0.A2 0.00338f
C1628 a_16458_15532# a_17800_15272# 0
C1629 sg13_inv_1_0.Y sg13_inv_1_1.Y 0.11018f
C1630 a_14859_16007# sg13_dfrbpq_1_3.Q 0
C1631 a_15856_16238# a_16266_15996# 0.10373f
C1632 sg13_inv_1_1.A sg13_dfrbpq_1_0.CLK 0.115f
C1633 sg13_dfrbpq_1_3.D a_14949_15213# 0.01365f
C1634 a_14506_15457# a_15051_15356# 0.01f
C1635 a_13499_15996# sg13_dfrbpq_1_4.D 0.15756f
C1636 sg13_nor2_1_0.A a_11595_16007# 0.00277f
C1637 a_12326_16746# a_12969_17137# 0.00801f
C1638 sg13_a21o_1_0.X VDD 0.97223f
C1639 sg13_a21oi_1_0.A1 a_14912_16878# 0.01629f
C1640 a_14340_15234# sg13_dfrbpq_1_0.CLK 0
C1641 sg13_a22oi_1_0.B2 a_15496_16878# 0.00165f
C1642 a_12335_16357# sg13_nor2_1_0.Y 0.02444f
C1643 a_14820_15247# a_15409_15255# 0
C1644 a_14340_16000# a_14314_15964# 0.36952f
C1645 sc_en clk_gating_en 4.07324f
C1646 a_16458_15532# a_16832_15366# 0.01061f
C1647 sg13_dfrbpq_1_3.D a_16048_15454# 0.00678f
C1648 a_14532_15552# a_15051_13844# 0
C1649 a_14949_15213# a_14949_13701# 0.00237f
C1650 sg13_nor2_1_0.A a_11953_15998# 0.00112f
C1651 a_15916_16119# sg13_inv_1_0.Y 0.01227f
C1652 sg13_dfrbpq_1_0.CLK a_12420_16746# 0
C1653 adc_en a_13576_4688# 0.24499f
C1654 a_13105_13799# sg13_a21o_1_0.X 0
C1655 sg13_a21oi_1_0.A1 a_11493_16007# 0
C1656 a_13131_16868# a_14128_16966# 0.02979f
C1657 a_12326_16746# a_12612_17064# 0.41329f
C1658 a_17696_15156# VDD 0
C1659 a_14820_15247# sg13_dfrbpq_1_0.CLK 0.00273f
C1660 a_13777_16823# a_13871_16823# 0.28931f
C1661 a_13838_12256# sg13_inv_1_0.Y 0
C1662 a_12900_16759# a_12326_16746# 0.31978f
C1663 a_14248_4688# VDD 0.25323f
C1664 sg13_a21o_1_0.A2 a_14155_12256# 0
C1665 a_14152_5498# Timer_en 0.00952f
C1666 a_16458_15532# sg13_dfrbpq_1_5.Q 0
C1667 a_14628_16421# a_14314_15964# 0.00463f
C1668 a_14859_16007# a_14054_16434# 0.097f
C1669 a_15791_15311# a_15051_13844# 0
C1670 a_15051_15356# a_15791_13799# 0
C1671 sg13_dfrbpq_1_3.D a_15409_15255# 0.0028f
C1672 sg13_nor2_1_0.A a_11940_14040# 0
C1673 sg13_a21oi_1_0.A1 a_13002_15996# 0
C1674 a_14757_16007# VDD 0.23714f
C1675 adc_en a_13960_4572# 0.00616f
C1676 adc_start a_25768_14914# 0
C1677 a_12708_14909# VDD 0.00957f
C1678 a_13131_16868# sg13_dfrbpq_1_0.CLK 0.0152f
C1679 a_14532_15552# sg13_nor2_1_0.B 0
C1680 a_14314_15964# sg13_a21oi_1_0.A2 0
C1681 sg13_nor2_1_0.A sg13_inv_1_0.Y 0.23317f
C1682 sg13_dfrbpq_1_3.D sg13_dfrbpq_1_0.CLK 0.08756f
C1683 a_8968_13760# VDD 0.25079f
C1684 a_14144_4572# VDD 0.00218f
C1685 a_13489_16767# sg13_dfrbpq_1_0.CLK 0.00932f
C1686 sg13_a21oi_1_0.A1 a_14538_17044# 0.14109f
C1687 a_16048_15454# a_16048_13942# 0
C1688 sg13_a21o_1_1.A2 a_17696_15366# 0
C1689 a_15217_16349# VDD 0.0014f
C1690 sg13_a22oi_1_0.B2 a_16735_16388# 0
C1691 sg13_dfrbpq_1_0.CLK a_10884_16434# 0
C1692 a_14144_23642# VDD 0.08585f
C1693 tx_start a_15688_25154# 0.00116f
C1694 a_15505_16357# sg13_inv_1_0.Y 0
C1695 sg13_dfrbpq_1_6.D a_12969_17137# 0
C1696 a_14098_14922# VDD 0
C1697 sg13_a22oi_1_0.B2 sg13_a21oi_1_0.A1 0.59937f
C1698 a_14949_13701# sg13_dfrbpq_1_0.CLK 0.27492f
C1699 a_12228_13735# sg13_buf_1_0.A 0
C1700 a_14949_15213# sg13_inv_1_0.Y 0.03847f
C1701 a_13499_15996# a_13601_16344# 0
C1702 a_13029_16725# a_13002_15996# 0.00351f
C1703 sg13_dfrbpq_1_0.CLK a_11595_16007# 0.03079f
C1704 a_10790_16434# a_11493_16007# 0.02432f
C1705 sg13_dfrbpq_1_3.D a_15409_14018# 0
C1706 sg13_dfrbpq_1_6.D a_12612_17064# 0.03855f
C1707 a_16048_13942# sg13_dfrbpq_1_0.CLK 0.00169f
C1708 a_13936_14726# a_13881_14607# 0.00412f
C1709 a_12939_14495# a_13996_14607# 0
C1710 a_12900_16759# sg13_dfrbpq_1_6.D 0.00768f
C1711 a_14188_17061# a_13131_16868# 0
C1712 sg13_o21ai_1_0.A1 a_12612_17064# 0
C1713 a_15993_15549# sg13_a22oi_1_0.B2 0
C1714 sg13_nor2b_1_0.Y a_12326_16746# 0
C1715 a_16048_15454# sg13_inv_1_0.Y 0.10177f
C1716 a_15599_16357# a_15784_14570# 0
C1717 a_11302_16421# a_11364_16421# 0
C1718 a_11493_16007# a_11953_16349# 0.02396f
C1719 a_11076_16000# a_11595_16007# 0.34102f
C1720 a_14859_16007# sg13_inv_1_1.Y 0
C1721 a_14949_13701# a_15409_14018# 0.01483f
C1722 a_13480_10830# sg13_a21o_1_0.X 0
C1723 sg13_dfrbpq_1_0.CLK a_11953_15998# 0
C1724 reset a_9728_13854# 0
C1725 sg13_inv_1_0.Y a_14128_16966# 0.10284f
C1726 sg13_buf_1_0.A a_13881_14607# 0
C1727 a_15409_13743# sg13_dfrbpq_1_0.CLK 0.00116f
C1728 sg13_dfrbpq_1_5.Q sg13_dfrbpq_1_6.D 0.02139f
C1729 a_15409_15255# sg13_inv_1_0.Y 0.00111f
C1730 sg13_nor2_1_0.A a_12134_14922# 0.002f
C1731 a_14152_10736# timer_done 0.26916f
C1732 a_14314_15964# VDD 0.11474f
C1733 sg13_dfrbpq_1_0.CLK a_11940_14040# 0.10394f
C1734 a_15051_13844# a_16108_14037# 0
C1735 sg13_dfrbpq_1_4.D a_13601_16344# 0.00663f
C1736 a_15856_16238# a_15801_16119# 0.00412f
C1737 a_14859_16007# a_15916_16119# 0
C1738 a_11595_16007# a_12335_16357# 0.26905f
C1739 wake_up_sg a_10024_15996# 0.26381f
C1740 a_11076_16000# a_11953_15998# 0
C1741 sg13_o21ai_1_0.A1 sg13_dfrbpq_1_5.Q 0.18261f
C1742 sg13_nor2_1_0.Y a_12394_14452# 0
C1743 a_15217_15998# sg13_o21ai_1_0.B1 0
C1744 sg13_inv_1_0.Y sg13_dfrbpq_1_0.CLK 0.58539f
C1745 a_15599_16357# a_15680_16878# 0
C1746 sg13_a21oi_1_0.A1 a_14437_17878# 0.00526f
C1747 a_12537_16119# sg13_nor2_1_0.A 0
C1748 adc_en VDD 0.14946f
C1749 a_12046_15276# a_11595_16007# 0
C1750 a_13702_12532# sg13_buf_1_0.A 0.09708f
C1751 sg13_dfrbpq_1_0.CLK a_13199_13799# 0.05264f
C1752 a_16048_13942# a_16458_14020# 0.10373f
C1753 a_15051_13844# a_15697_13799# 0.00647f
C1754 a_14440_5412# timer_done 0.05144f
C1755 a_12592_16238# sg13_nor2_1_0.B 0
C1756 a_12241_16357# a_12754_16434# 0
C1757 a_13499_15996# sg13_nor2_1_0.Y 0.00414f
C1758 a_14506_13945# a_14246_13722# 0.75507f
C1759 a_14440_5412# a_14632_4688# 0
C1760 a_14152_5498# a_14248_4688# 0
C1761 sg13_dfrbpq_1_6.D a_12754_16434# 0
C1762 sg13_inv_1_0.Y a_11076_16000# 0.38728f
C1763 sg13_a21oi_1_0.A1 a_12420_14488# 0
C1764 sg13_buf_1_4.A VDD 0.91842f
C1765 sg13_nor2b_1_0.Y a_12241_16357# 0
C1766 sg13_inv_1_1.A a_16430_14832# 0
C1767 a_15051_15356# a_14757_16007# 0
C1768 a_15409_14018# sg13_inv_1_0.Y 0.01621f
C1769 sg13_nor2b_1_0.Y sg13_dfrbpq_1_6.D 0.00172f
C1770 a_14859_16007# a_15505_16357# 0.00647f
C1771 sg13_inv_1_0.Y a_12335_16357# 0.16804f
C1772 a_12268_15532# sg13_nor2b_1_0.Y 0.01673f
C1773 sg13_inv_1_1.A a_13936_14726# 0.00238f
C1774 sg13_a21oi_1_0.A1 a_13864_16082# 0.00342f
C1775 adc_start sg13_dfrbpq_1_1.Q 0.008f
C1776 sg13_a21o_1_1.A2 VDD 0.50225f
C1777 sg13_a21oi_1_0.A1 a_13679_14845# 0
C1778 a_13866_14020# sg13_inv_1_1.Y 0
C1779 uart_busy a_15976_25068# 0.26742f
C1780 a_10024_15996# sg13_dfrbpq_1_4.D 0.00179f
C1781 a_14152_5842# sg13_buf_1_0.A 0.00233f
C1782 sg13_nor2_1_0.B a_12357_13701# 0.00142f
C1783 a_14532_15552# a_15856_16238# 0
C1784 a_14949_15213# a_14859_16007# 0.00237f
C1785 a_16458_14020# sg13_inv_1_0.Y 0
C1786 a_14188_17061# sg13_inv_1_0.Y 0.01227f
C1787 a_14506_13945# a_14820_13735# 0.00463f
C1788 a_14246_15234# sg13_buf_1_0.A 0
C1789 sg13_a22oi_1_0.B2 a_15976_25068# 0.24834f
C1790 a_14144_23986# sg13_a21oi_1_0.A2 0.00131f
C1791 sg13_dfrbpq_1_4.D sg13_nor2_1_0.Y 0.22754f
C1792 a_15599_16357# sg13_inv_1_1.A 0.00294f
C1793 a_12046_15276# sg13_inv_1_0.Y 0.00348f
C1794 sg13_buf_1_0.A a_14336_5498# 0.02549f
C1795 sg13_inv_1_1.A sg13_buf_1_0.A 0.00165f
C1796 sg13_a21oi_1_0.A1 a_14235_17564# 0.27988f
C1797 sg13_nor2b_1_0.Y a_12297_14113# 0
C1798 sg13_a21oi_1_0.A1 a_16266_15996# 0
C1799 a_11654_13722# a_12817_14018# 0
C1800 a_11940_14040# a_12459_13844# 0.34114f
C1801 a_14998_16742# VDD 0.01065f
C1802 a_15791_15311# a_15856_16238# 0
C1803 sg13_dfrbpq_1_0.CLK a_12134_14922# 0.00446f
C1804 sg13_inv_1_0.Y a_12459_13844# 0.48314f
C1805 sg13_dfrbpq_1_5.Q sg13_o21ai_1_0.B1 0.00279f
C1806 sg13_dfrbpq_1_1.Q a_16051_14746# 0.22317f
C1807 a_14506_13945# sg13_and2_1_0.X 0.00937f
C1808 a_12357_13701# a_13456_13942# 0
C1809 a_12459_13844# a_13199_13799# 0.26905f
C1810 a_12537_16119# sg13_dfrbpq_1_0.CLK 0
C1811 a_13864_16082# a_13029_16725# 0.00104f
C1812 a_25672_11890# VDD 0.00121f
C1813 a_25856_16668# VDD 0
C1814 sg13_dfrbpq_1_0.CLK a_13297_14837# 0.00575f
C1815 a_14757_16007# a_14912_16878# 0.00112f
C1816 a_15217_15998# a_14054_16434# 0
C1817 sg13_inv_1_0.Y a_13516_14037# 0.01414f
C1818 a_14155_12256# sg13_buf_1_4.A 0.00395f
C1819 sg13_dfrbpq_1_3.D a_13936_14726# 0
C1820 a_12326_16746# sg13_a21oi_1_0.A2 0.00214f
C1821 a_13199_13799# a_13516_14037# 0.00247f
C1822 a_14859_16007# sg13_dfrbpq_1_0.CLK 0.0562f
C1823 sg13_dfrbpq_1_0.CLK a_12777_14531# 0
C1824 a_12335_16357# a_12134_14922# 0
C1825 a_14073_17061# sg13_a21oi_1_0.A2 0.00165f
C1826 a_13664_10830# VDD 0.06411f
C1827 a_11914_13945# a_11654_13722# 0.75507f
C1828 a_16735_15972# sg13_a21o_1_1.A2 0.00131f
C1829 wake_up_sg a_11595_16007# 0
C1830 a_16832_15366# sg13_dfrbpq_1_3.Q 0.01342f
C1831 sg13_dfrbpq_1_3.D a_15599_16357# 0
C1832 a_14246_13722# a_14346_14484# 0
C1833 sg13_dfrbpq_1_3.D sg13_buf_1_0.A 0.00454f
C1834 sg13_inv_1_0.Y a_9728_13854# 0.00154f
C1835 a_14697_16043# VDD 0
C1836 a_13480_10830# sg13_buf_1_4.A 0.00195f
C1837 a_12046_15276# a_12134_14922# 0
C1838 a_12652_16119# a_12592_16238# 0.01042f
C1839 a_12537_16119# a_12335_16357# 0.00689f
C1840 a_13131_16868# sg13_dfrbpq_1_4.D 0
C1841 Timer_en a_13960_4782# 0.01683f
C1842 a_14144_23986# VDD 0.00293f
C1843 a_14340_16000# sg13_dfrbpq_1_6.D 0.0053f
C1844 sg13_dfrbpq_1_3.Q sg13_dfrbpq_1_5.Q 0.46867f
C1845 sg13_inv_2_1.A a_17696_15156# 0
C1846 a_15409_15530# VDD 0.0077f
C1847 a_14144_17594# sg13_inv_1_0.Y 0
C1848 a_14061_12256# a_13838_12256# 0
C1849 a_14340_16000# sg13_o21ai_1_0.A1 0.00316f
C1850 a_12652_16119# sg13_nor2_1_0.B 0
C1851 sg13_nor2_1_0.B a_12939_14495# 0.00444f
C1852 sg13_a22oi_1_0.B2 a_14757_16007# 0.04061f
C1853 a_14628_16421# sg13_dfrbpq_1_6.D 0.0029f
C1854 a_16458_15532# VDD 0.38282f
C1855 sg13_inv_1_0.Y a_12394_14452# 0.27901f
C1856 a_14061_12256# a_14152_10736# 0
C1857 sg13_inv_1_1.A a_15784_14570# 0
C1858 wake_up_sg sg13_inv_1_0.Y 0.00145f
C1859 a_12357_13701# a_12939_14495# 0
C1860 sg13_a21oi_1_0.A1 a_13864_16426# 0.00382f
C1861 sg13_dfrbpq_1_4.D a_11595_16007# 0.02579f
C1862 sg13_nor2_1_0.B a_13297_14486# 0
C1863 sg13_dfrbpq_1_6.D sg13_a21oi_1_0.A2 0.05283f
C1864 a_12326_16746# VDD 0.7807f
C1865 sg13_a22oi_1_0.B2 a_15217_16349# 0.00677f
C1866 a_16210_15234# VDD 0
C1867 sg13_o21ai_1_0.A1 sg13_a21oi_1_0.A2 0
C1868 a_11914_13945# sg13_a21o_1_0.X 0.00113f
C1869 a_14073_17061# VDD 0.00274f
C1870 sg13_inv_1_0.Y a_13936_14726# 0.10353f
C1871 a_15791_15311# a_16051_14746# 0
C1872 a_11940_14040# sg13_buf_1_0.A 0.00175f
C1873 a_13866_14020# sg13_dfrbpq_1_0.CLK 0.00307f
C1874 a_13199_13799# a_13936_14726# 0
C1875 a_13456_13942# a_12939_14495# 0
C1876 sg13_and2_1_0.X a_14346_14484# 0
C1877 sg13_dfrbpq_1_4.D a_11953_15998# 0.00363f
C1878 a_15599_16357# sg13_inv_1_0.Y 0.13423f
C1879 a_15096_17064# VDD 0.01832f
C1880 sg13_inv_1_0.Y sg13_buf_1_0.A 0.69243f
C1881 a_13768_10736# a_13664_10620# 0
C1882 a_13480_10830# a_13664_10830# 0.0524f
C1883 a_13199_13799# sg13_buf_1_0.A 0.0145f
C1884 adc_start a_15051_13844# 0
C1885 a_15697_15311# sg13_a21o_1_1.A2 0
C1886 a_11302_16421# VDD 0
C1887 sg13_dfrbpq_1_6.D a_14148_16434# 0
C1888 a_12612_17064# sg13_inv_1_1.Y 0
C1889 a_14538_17044# a_14314_15964# 0
C1890 sg13_dfrbpq_1_3.D a_15784_14570# 0.02888f
C1891 sg13_dfrbpq_1_0.CLK a_15784_14914# 0.00347f
C1892 sg13_inv_1_0.Y sg13_dfrbpq_1_4.D 0.15656f
C1893 a_13618_13722# VDD 0
C1894 sg13_buf_1_6.X a_9728_13854# 0.02132f
C1895 a_14340_16000# sg13_o21ai_1_0.B1 0
C1896 clk_gating_en VDD 0.20604f
C1897 a_14440_5412# sc_en 0.24441f
C1898 a_12134_14922# a_12394_14452# 0.75507f
C1899 a_12241_16357# VDD 0
C1900 sg13_inv_1_1.A sg13_nor2_1_0.Y 0
C1901 sg13_a22oi_1_0.B2 a_14314_15964# 0.00142f
C1902 a_13105_13799# a_13618_13722# 0
C1903 adc_done adc_start 0.00514f
C1904 sg13_dfrbpq_1_6.D VDD 0.58292f
C1905 a_14532_14040# sg13_dfrbpq_1_1.Q 0
C1906 a_14949_13701# a_15784_14570# 0.00171f
C1907 a_15993_14037# VDD 0
C1908 a_14628_16421# sg13_o21ai_1_0.B1 0
C1909 a_12268_15532# VDD 0.00713f
C1910 a_14912_16668# sg13_dfrbpq_1_0.CLK 0
C1911 sg13_o21ai_1_0.A1 VDD 0.45976f
C1912 a_14248_4688# a_13960_4782# 0.00536f
C1913 a_14246_15234# sg13_inv_1_1.A 0.02125f
C1914 a_12420_14488# a_12708_14909# 0.43707f
C1915 a_14248_23556# tx_start 0.2541f
C1916 a_14532_15552# sg13_a21oi_1_0.A1 0
C1917 adc_start a_15697_13799# 0
C1918 a_15688_25498# VDD 0.00207f
C1919 a_16210_13722# sg13_and2_1_0.X 0
C1920 a_14912_16878# a_14998_16742# 0
C1921 sg13_o21ai_1_0.B1 sg13_a21oi_1_0.A2 0.0284f
C1922 a_14246_15234# a_14340_15234# 0.00716f
C1923 a_15051_15356# a_15409_15530# 0.02138f
C1924 a_14340_16000# a_14566_16421# 0.0052f
C1925 a_15791_13799# sg13_dfrbpq_1_1.Q 0.0075f
C1926 a_12228_13735# a_11940_14040# 0.43707f
C1927 a_25856_17938# VDD 0
C1928 a_17024_13644# VDD 0
C1929 a_14506_13945# VDD 0.10142f
C1930 a_7816_15996# sg13_dfrbpq_1_0.CLK 0.2561f
C1931 a_12394_14452# a_12777_14531# 0.00333f
C1932 a_12837_14495# a_13585_14845# 0.01058f
C1933 sg13_nor2_1_0.A a_12612_17064# 0
C1934 a_12297_14113# VDD 0
C1935 timer_done sg13_buf_1_0.A 0.34877f
C1936 a_12228_13735# sg13_inv_1_0.Y 0.01622f
C1937 a_17128_13760# sg13_a21o_1_1.A2 0
C1938 sg13_dfrbpq_1_5.Q a_15680_16668# 0.0013f
C1939 sg13_buf_1_0.A a_14632_4688# 0.24846f
C1940 a_12650_15532# sg13_nor2_1_0.A 0
C1941 a_13401_14037# a_13456_13942# 0.00412f
C1942 a_13131_16868# sg13_nor2_1_0.Y 0.00365f
C1943 a_14246_15234# a_14820_15247# 0.31978f
C1944 a_14340_16000# sg13_dfrbpq_1_3.Q 0
C1945 a_14566_16421# a_14628_16421# 0
C1946 sg13_a21oi_1_0.A1 a_13871_16823# 0.01324f
C1947 uart_done sg13_a21oi_1_0.A2 0.03225f
C1948 a_14820_15247# sg13_inv_1_1.A 0.0019f
C1949 sg13_inv_2_1.A sg13_a21o_1_1.A2 0.23726f
C1950 sg13_dfrbpq_1_3.D sg13_nor2_1_0.Y 0
C1951 a_13679_14845# a_14098_14922# 0.00174f
C1952 a_12939_14495# a_13297_14486# 0.02138f
C1953 sg13_a22oi_1_0.B2 sg13_a21o_1_1.A2 0
C1954 a_14758_15247# sg13_a21oi_1_0.A1 0
C1955 sg13_buf_1_5.X a_13768_10736# 0.00702f
C1956 a_14144_23642# a_13960_25068# 0
C1957 a_14566_16421# sg13_a21oi_1_0.A2 0
C1958 a_16840_13644# sg13_a21o_1_1.A2 0
C1959 a_15791_15311# a_15993_15549# 0.00689f
C1960 a_14859_16007# a_15599_16357# 0.26905f
C1961 a_14538_17044# a_14998_16742# 0
C1962 sg13_inv_1_0.Y a_15784_14570# 0
C1963 a_15217_15998# sg13_dfrbpq_1_0.CLK 0.00669f
C1964 sg13_inv_1_1.A a_13131_16868# 0
C1965 a_14506_15457# a_14532_15552# 0.36952f
C1966 sg13_dfrbpq_1_3.D a_14246_15234# 0.28605f
C1967 a_12537_16119# sg13_dfrbpq_1_4.D 0.00153f
C1968 sg13_dfrbpq_1_4.D a_13297_14837# 0
C1969 sg13_dfrbpq_1_3.D sg13_inv_1_1.A 0.49583f
C1970 sg13_inv_1_0.Y a_13881_14607# 0.00451f
C1971 a_15505_16357# sg13_dfrbpq_1_5.Q 0.00389f
C1972 sg13_a22oi_1_0.B2 a_14998_16742# 0.10281f
C1973 sg13_a21oi_1_0.A1 a_13777_16823# 0.00351f
C1974 a_13856_25154# sg13_a21oi_1_0.A2 0
C1975 a_9728_13644# VDD 0
C1976 a_14889_15625# sg13_dfrbpq_1_0.CLK 0
C1977 a_13768_10736# Timer_en 0.24441f
C1978 a_11595_16007# sg13_nor2_1_0.Y 0
C1979 a_14340_16000# a_14054_16434# 0.41329f
C1980 a_14949_15213# sg13_dfrbpq_1_5.Q 0
C1981 sg13_dfrbpq_1_3.D a_14340_15234# 0
C1982 a_14859_16007# sg13_dfrbpq_1_4.D 0
C1983 a_12166_13735# sg13_a21o_1_0.X 0
C1984 sg13_o21ai_1_0.B1 VDD 0.6707f
C1985 a_13029_16725# a_13871_16823# 0.00332f
C1986 a_12612_17064# a_14128_16966# 0.00242f
C1987 a_16832_15156# VDD 0
C1988 a_13702_12532# sg13_inv_1_0.Y 0
C1989 a_14336_5842# Timer_en 0
C1990 a_13459_12404# a_13838_12256# 0
C1991 a_15697_15311# a_16210_15234# 0
C1992 a_14628_16421# a_14054_16434# 0.31978f
C1993 sg13_nor2b_1_0.Y sg13_nor2_1_0.A 0.22641f
C1994 sg13_dfrbpq_1_3.D a_14820_15247# 0.00833f
C1995 adc_en a_13960_4782# 0.02118f
C1996 sg13_a21oi_1_0.A1 a_12592_16238# 0
C1997 a_14314_15964# a_13679_14845# 0
C1998 a_12837_14495# VDD 0.26539f
C1999 a_13029_16725# a_13489_17042# 0.01483f
C2000 a_12612_17064# sg13_dfrbpq_1_0.CLK 0.0952f
C2001 sg13_inv_1_1.A a_16048_13942# 0
C2002 a_16832_15366# sg13_dfrbpq_1_0.CLK 0
C2003 a_10024_15996# sg13_inv_1_0.Y 0
C2004 uart_done VDD 0.20954f
C2005 a_13489_16767# a_13131_16868# 0.00104f
C2006 a_12900_16759# sg13_dfrbpq_1_0.CLK 0.00481f
C2007 a_13777_16823# a_13029_16725# 0.01058f
C2008 a_16294_14484# VDD 0.37801f
C2009 a_14054_16434# sg13_a21oi_1_0.A2 0.00243f
C2010 a_14144_4782# VDD 0.06713f
C2011 a_13866_14020# a_13936_14726# 0
C2012 a_13105_13799# a_12837_14495# 0
C2013 a_15791_15311# a_15791_13799# 0
C2014 sg13_inv_1_0.Y sg13_nor2_1_0.Y 0.75458f
C2015 sg13_a21oi_1_0.A1 sg13_nor2_1_0.B 0
C2016 a_15051_15356# sg13_o21ai_1_0.A1 0
C2017 a_14566_16421# VDD 0
C2018 a_12326_16746# a_11493_16007# 0
C2019 a_14346_14484# VDD 0.40857f
C2020 tx_start a_15872_25498# 0
C2021 a_14246_13722# sg13_dfrbpq_1_0.CLK 0.00363f
C2022 sg13_dfrbpq_1_5.Q sg13_dfrbpq_1_0.CLK 0.00304f
C2023 a_15409_15530# sg13_a22oi_1_0.B2 0.00156f
C2024 a_14246_15234# sg13_inv_1_0.Y 0.11855f
C2025 a_13866_14020# sg13_buf_1_0.A 0.05756f
C2026 sg13_buf_1_4.A a_13679_14845# 0
C2027 a_13856_25154# VDD 0.09174f
C2028 reset sg13_inv_1_0.Y 0
C2029 a_16840_13854# sg13_a21o_1_1.A2 0.0012f
C2030 sg13_dfrbpq_1_3.Q VDD 0.64661f
C2031 a_14340_16000# sg13_inv_1_1.Y 0.00528f
C2032 a_10790_16434# a_11050_15964# 0.75507f
C2033 a_13192_12132# sg13_a21o_1_0.X 0.00379f
C2034 sg13_dfrbpq_1_3.D a_14949_13701# 0.00226f
C2035 sg13_dfrbpq_1_0.CLK a_11364_16421# 0.00868f
C2036 a_12612_17064# a_12335_16357# 0.00248f
C2037 sg13_inv_1_1.A sg13_inv_1_0.Y 0.07242f
C2038 a_12136_16878# a_12326_16746# 0.00201f
C2039 a_12900_16759# a_12335_16357# 0
C2040 a_16458_15532# sg13_inv_2_1.A 0.00627f
C2041 a_16458_15532# sg13_a22oi_1_0.B2 0.00158f
C2042 a_14054_16434# a_14148_16434# 0.00716f
C2043 a_14340_15234# sg13_inv_1_0.Y 0
C2044 a_14246_13722# a_15409_14018# 0
C2045 a_14532_14040# a_15051_13844# 0.34114f
C2046 a_15697_15311# sg13_o21ai_1_0.A1 0
C2047 a_14628_16421# sg13_inv_1_1.Y 0
C2048 sg13_nor2_1_0.A a_11464_13854# 0
C2049 sg13_dfrbpq_1_0.CLK a_12754_16434# 0
C2050 a_11076_16000# a_11364_16421# 0.43707f
C2051 sg13_dfrbpq_1_3.D a_16048_13942# 0
C2052 a_13029_16725# sg13_nor2_1_0.B 0.00197f
C2053 a_15856_16238# a_16051_14746# 0
C2054 reset a_8776_13854# 0.03394f
C2055 sg13_inv_1_0.Y a_12420_16746# 0
C2056 a_14820_13735# sg13_dfrbpq_1_0.CLK 0
C2057 a_14506_15457# sg13_nor2_1_0.B 0
C2058 uart_done a_13856_25498# 0.00127f
C2059 sg13_inv_1_1.Y sg13_a21oi_1_0.A2 0.02467f
C2060 a_14912_16878# sg13_dfrbpq_1_6.D 0.0023f
C2061 a_14820_15247# sg13_inv_1_0.Y 0.00549f
C2062 a_14054_16434# VDD 0.80787f
C2063 sg13_nor2b_1_0.Y sg13_dfrbpq_1_0.CLK 0
C2064 sg13_dfrbpq_1_3.D a_15409_13743# 0
C2065 wake_up_sg a_7816_15996# 0.01128f
C2066 a_11050_15964# a_11433_16043# 0.00333f
C2067 a_14949_13701# a_16048_13942# 0
C2068 a_15051_13844# a_15791_13799# 0.26905f
C2069 a_11493_16007# a_12241_16357# 0.01058f
C2070 sg13_o21ai_1_0.A1 a_14912_16878# 0.02686f
C2071 sg13_dfrbpq_1_6.D a_11493_16007# 0.00154f
C2072 sg13_nor2_1_0.Y a_12134_14922# 0
C2073 a_14859_16007# a_15680_16878# 0.00105f
C2074 a_16210_13722# VDD 0
C2075 sg13_inv_1_0.Y a_13131_16868# 0.42194f
C2076 a_13459_12404# sg13_dfrbpq_1_0.CLK 0
C2077 a_14061_12256# sg13_buf_1_0.A 0
C2078 sg13_nor2b_1_0.Y a_11076_16000# 0.00296f
C2079 a_13489_16767# sg13_inv_1_0.Y 0
C2080 sg13_and2_1_0.X sg13_dfrbpq_1_0.CLK 0
C2081 sg13_a22oi_1_0.B2 a_15096_17064# 0.01073f
C2082 a_14152_5842# timer_done 0.00274f
C2083 a_12335_16357# a_12754_16434# 0.00174f
C2084 sg13_dfrbpq_1_3.Q a_16735_15972# 0.02037f
C2085 sg13_dfrbpq_1_3.D sg13_inv_1_0.Y 0.12721f
C2086 a_15051_15356# sg13_o21ai_1_0.B1 0
C2087 a_11595_16007# a_11953_15998# 0.02138f
C2088 a_15791_13799# a_16108_14037# 0.00247f
C2089 a_14532_14040# a_15697_13799# 0.43239f
C2090 a_14949_13701# a_15409_13743# 0.02396f
C2091 sg13_dfrbpq_1_6.D a_13002_15996# 0.00209f
C2092 a_14340_16000# a_15505_16357# 0.43239f
C2093 sg13_nor2_1_0.Y a_13297_14837# 0
C2094 timer_done a_14336_5498# 0.00114f
C2095 a_12136_16878# sg13_dfrbpq_1_6.D 0.03359f
C2096 a_12817_13743# VDD 0.0013f
C2097 sg13_nor2b_1_0.Y a_12335_16357# 0
C2098 a_14949_13701# sg13_inv_1_0.Y 0.03758f
C2099 a_14532_15552# a_14757_16007# 0
C2100 a_14949_15213# a_14340_16000# 0
C2101 a_14538_17044# sg13_dfrbpq_1_6.D 0.01463f
C2102 a_15791_13799# a_15697_13799# 0.28931f
C2103 a_14506_13945# a_14889_14113# 0.00333f
C2104 a_14152_5498# a_14144_4782# 0
C2105 a_14538_17044# sg13_o21ai_1_0.A1 0.00167f
C2106 a_12046_15276# sg13_nor2b_1_0.Y 0.30331f
C2107 sg13_inv_1_0.Y a_11595_16007# 0.4356f
C2108 reset sg13_buf_1_6.X 0.00507f
C2109 sg13_a22oi_1_0.B2 sg13_dfrbpq_1_6.D 0.10701f
C2110 uart_busy a_15688_25498# 0.00347f
C2111 sg13_nor2_1_0.B a_11654_13722# 0
C2112 a_13480_10620# sg13_buf_1_0.A 0.00274f
C2113 a_16048_13942# sg13_inv_1_0.Y 0.10167f
C2114 sc_en sg13_buf_1_0.A 0.17176f
C2115 sg13_inv_1_1.Y VDD 0.58576f
C2116 a_17024_13644# a_17128_13760# 0
C2117 sg13_a22oi_1_0.B2 sg13_o21ai_1_0.A1 0.28907f
C2118 a_14859_16007# sg13_inv_1_1.A 0.00517f
C2119 sg13_a22oi_1_0.B2 a_15688_25498# 0
C2120 sg13_a21oi_1_0.A1 a_15856_16238# 0
C2121 a_11654_13722# a_12357_13701# 0.02454f
C2122 sg13_inv_1_0.Y a_11953_15998# 0.01783f
C2123 tx_start sg13_a21oi_1_0.A2 0.10845f
C2124 a_15976_25068# a_15872_25154# 0.00624f
C2125 a_14912_16878# sg13_o21ai_1_0.B1 0
C2126 a_15916_16119# VDD 0.00728f
C2127 sg13_inv_1_0.Y a_11940_14040# 0.41511f
C2128 a_11940_14040# a_13199_13799# 0.01529f
C2129 sg13_dfrbpq_1_1.Q sg13_a21o_1_1.A2 0.01021f
C2130 a_15680_16668# VDD 0
C2131 a_14340_16000# sg13_dfrbpq_1_0.CLK 0.11238f
C2132 a_13838_12256# VDD 0
C2133 a_16108_15549# sg13_dfrbpq_1_3.Q 0
C2134 a_16458_15532# a_16266_15996# 0
C2135 sg13_inv_1_0.Y a_13199_13799# 0.15132f
C2136 a_14128_16966# sg13_a21oi_1_0.A2 0.0045f
C2137 a_14628_16421# sg13_dfrbpq_1_0.CLK 0.00448f
C2138 a_12652_16119# a_10790_16434# 0
C2139 a_14152_10736# VDD 0.24333f
C2140 sg13_nor2_1_0.A VDD 0.89006f
C2141 a_15697_15311# sg13_dfrbpq_1_3.Q 0
C2142 sg13_dfrbpq_1_0.CLK a_13585_14845# 0.00879f
C2143 a_14437_17878# sg13_dfrbpq_1_6.D 0
C2144 a_13768_10736# sg13_buf_1_4.A 0.26372f
C2145 a_14538_17044# sg13_o21ai_1_0.B1 0.00196f
C2146 sg13_inv_1_0.Y a_8776_13854# 0
C2147 sg13_dfrbpq_1_0.CLK sg13_a21oi_1_0.A2 0.21854f
C2148 a_15505_16357# VDD 0.00179f
C2149 a_12537_16119# a_11595_16007# 0
C2150 a_25768_25498# VDD 0.00121f
C2151 Timer_en a_13472_4782# 0
C2152 a_14290_16746# sg13_a21oi_1_0.A2 0
C2153 a_12612_17064# sg13_dfrbpq_1_4.D 0
C2154 a_11914_13945# a_12297_14113# 0.00333f
C2155 sg13_a21o_1_0.X a_12357_13701# 0.00165f
C2156 a_14440_5412# VDD 0.26621f
C2157 sg13_a22oi_1_0.B2 sg13_o21ai_1_0.B1 0.84375f
C2158 sg13_inv_1_1.A a_13866_14020# 0
C2159 a_15599_16357# sg13_dfrbpq_1_5.Q 0.00807f
C2160 tx_start VDD 0.71931f
C2161 a_14949_15213# VDD 0.25572f
C2162 a_12650_15532# sg13_dfrbpq_1_4.D 0
C2163 a_14246_13722# sg13_buf_1_0.A 0.03879f
C2164 a_14061_12256# a_13702_12532# 0.01325f
C2165 sg13_nor2b_1_0.Y a_12394_14452# 0
C2166 a_13871_16823# a_14314_15964# 0
C2167 sg13_a21o_1_0.X a_13456_13942# 0
C2168 sg13_nor2_1_0.B a_12708_14909# 0.00303f
C2169 a_13864_16082# sg13_dfrbpq_1_6.D 0
C2170 a_16048_15454# VDD 0.16077f
C2171 a_14340_13722# sg13_buf_1_0.A 0
C2172 sg13_inv_1_0.Y a_12134_14922# 0.1319f
C2173 a_14128_16966# VDD 0.18514f
C2174 sg13_dfrbpq_1_4.D a_11364_16421# 0
C2175 a_12537_16119# sg13_inv_1_0.Y 0.0058f
C2176 a_14188_17061# sg13_a21oi_1_0.A2 0.00197f
C2177 a_14235_17564# sg13_dfrbpq_1_6.D 0.00109f
C2178 a_15409_15255# VDD 0.00121f
C2179 sg13_inv_1_0.Y a_13297_14837# 0.00217f
C2180 sg13_and2_1_0.X a_13936_14726# 0
C2181 a_15791_15311# sg13_a21o_1_1.A2 0.00424f
C2182 sg13_inv_1_0.Y sg13_buf_1_6.X 0.12144f
C2183 sg13_dfrbpq_1_3.Q sg13_inv_2_1.A 0.11219f
C2184 sg13_dfrbpq_1_0.CLK VDD 1.90753f
C2185 sg13_a22oi_1_0.B2 sg13_dfrbpq_1_3.Q 0.14335f
C2186 a_16458_15532# sg13_dfrbpq_1_1.Q 0.00135f
C2187 a_14859_16007# sg13_inv_1_0.Y 0.426f
C2188 a_14290_16746# VDD 0.00129f
C2189 sg13_inv_1_0.Y a_12777_14531# 0
C2190 a_13768_10736# a_13664_10830# 0.00624f
C2191 a_14437_17878# sg13_o21ai_1_0.B1 0.00593f
C2192 a_13459_12404# sg13_buf_1_0.A 0.23676f
C2193 a_13105_13799# sg13_dfrbpq_1_0.CLK 0.01254f
C2194 sg13_nor2b_1_0.Y sg13_dfrbpq_1_4.D 0.00483f
C2195 sg13_and2_1_0.X sg13_buf_1_0.A 0.34242f
C2196 a_11076_16000# VDD 0.07813f
C2197 adc_start a_14532_14040# 0
C2198 sg13_buf_1_6.X a_8776_13854# 0
C2199 a_8968_13760# a_8776_13644# 0
C2200 a_15409_14018# VDD 0.00775f
C2201 a_14538_17044# a_14054_16434# 0
C2202 sg13_dfrbpq_1_3.D a_15784_14914# 0.00732f
C2203 adc_start a_15791_13799# 0
C2204 a_15505_16357# a_16018_16434# 0
C2205 a_12335_16357# VDD 0.17199f
C2206 sg13_a22oi_1_0.B2 a_14054_16434# 0.00267f
C2207 timer_done a_14632_4688# 0.02458f
C2208 a_16458_14020# VDD 0.38571f
C2209 a_14440_5412# a_14152_5498# 0.00524f
C2210 a_13576_4688# a_13472_4572# 0
C2211 a_14188_17061# VDD 0.01393f
C2212 a_12420_14488# a_12837_14495# 0.37583f
C2213 a_12046_15276# VDD 0.21597f
C2214 a_15217_15998# sg13_inv_1_1.A 0.00186f
C2215 a_12969_17137# sg13_nor2_1_0.Y 0
C2216 a_14949_15213# a_15051_15356# 0.47622f
C2217 a_14144_17594# sg13_a21oi_1_0.A2 0.02323f
C2218 a_14532_15552# a_15409_15530# 0
C2219 a_14246_15234# a_14889_15625# 0.00801f
C2220 power_on VSS 0.06665f
C2221 clk_gating_en VSS 1.21618f
C2222 uart_en VSS 0.70739f
C2223 adc_en VSS 1.23599f
C2224 sc_en VSS 0.67035f
C2225 Timer_en VSS 1.20789f
C2226 timer_done VSS 2.12396f
C2227 adc_start VSS 4.4762f
C2228 reset VSS 2.58111f
C2229 adc_done VSS 3.38427f
C2230 wake_up_sg VSS 1.88149f
C2231 clk VSS 2.61586f
C2232 tx_start VSS 1.6554f
C2233 uart_busy VSS 1.76724f
C2234 uart_done VSS 1.51195f
C2235 VDD VSS 1.38739p
C2236 a_25768_4572# VSS 0.02451f $ **FLOATING
C2237 a_25768_4782# VSS 0.1466f $ **FLOATING
C2238 a_14144_4572# VSS 0.00582f $ **FLOATING
C2239 a_13960_4572# VSS 0.01837f $ **FLOATING
C2240 a_14144_4782# VSS 0.03789f $ **FLOATING
C2241 a_13960_4782# VSS 0.08475f $ **FLOATING
C2242 a_13472_4572# VSS 0.00918f $ **FLOATING
C2243 a_13472_4782# VSS 0.06097f $ **FLOATING
C2244 a_14632_4688# VSS 0.36578f
C2245 a_14248_4688# VSS 0.36097f
C2246 a_13576_4688# VSS 0.3804f
C2247 a_14336_5498# VSS 0.03748f $ **FLOATING
C2248 a_14152_5498# VSS 0.09803f $ **FLOATING
C2249 a_14440_5412# VSS 0.37955f
C2250 a_14336_5842# VSS 0.00677f $ **FLOATING
C2251 a_14152_5842# VSS 0.02583f $ **FLOATING
C2252 a_13664_10620# VSS 0.00677f $ **FLOATING
C2253 a_13480_10620# VSS 0.02583f $ **FLOATING
C2254 a_13664_10830# VSS 0.03807f $ **FLOATING
C2255 a_13480_10830# VSS 0.09895f $ **FLOATING
C2256 a_14152_10736# VSS 0.36228f
C2257 a_13768_10736# VSS 0.36904f
C2258 a_25856_11546# VSS 0.07765f $ **FLOATING
C2259 a_25672_11546# VSS 0.09948f $ **FLOATING
C2260 a_25856_11890# VSS 0.00533f $ **FLOATING
C2261 a_25672_11890# VSS 0.02391f $ **FLOATING
C2262 a_14155_12256# VSS 0.00659f
C2263 a_13838_12256# VSS 0.01083f
C2264 a_13192_12132# VSS 0.02473f $ **FLOATING
C2265 a_13702_12532# VSS 0.02782f
C2266 a_13192_12342# VSS 0.09162f $ **FLOATING
C2267 a_14061_12256# VSS 0.30041f
C2268 sg13_buf_1_5.X VSS 1.23387f
C2269 sg13_a21o_1_0.A2 VSS 0.9063f
C2270 a_13459_12404# VSS 0.51073f
C2271 a_17024_13644# VSS 0.00585f $ **FLOATING
C2272 a_16840_13644# VSS 0.01821f $ **FLOATING
C2273 a_17024_13854# VSS 0.03753f $ **FLOATING
C2274 a_16840_13854# VSS 0.07982f $ **FLOATING
C2275 a_16210_13722# VSS 0.00329f
C2276 a_15697_13799# VSS 0.09498f
C2277 a_15409_13743# VSS 0.00443f
C2278 a_14820_13735# VSS 0.03599f
C2279 a_17128_13760# VSS 0.36807f
C2280 a_16458_14020# VSS 0.41792f
C2281 a_16048_13942# VSS 0.24416f
C2282 a_15791_13799# VSS 0.51893f
C2283 a_14340_13722# VSS 0
C2284 a_13618_13722# VSS 0.00329f
C2285 a_15051_13844# VSS 0.3698f
C2286 a_14949_13701# VSS 0.77467f
C2287 a_14532_14040# VSS 1.57593f
C2288 a_14246_13722# VSS 0.17149f
C2289 sg13_and2_1_0.X VSS 0.72237f
C2290 a_14506_13945# VSS 0.23698f
C2291 sg13_buf_1_4.A VSS 1.36477f
C2292 a_13105_13799# VSS 0.09495f
C2293 a_12817_13743# VSS 0.00443f
C2294 a_12228_13735# VSS 0.03599f
C2295 a_13866_14020# VSS 0.42028f
C2296 a_13456_13942# VSS 0.24478f
C2297 a_13199_13799# VSS 0.51866f
C2298 a_11748_13722# VSS 0
C2299 a_11464_13644# VSS 0.02444f $ **FLOATING
C2300 a_12459_13844# VSS 0.37091f
C2301 a_12357_13701# VSS 0.77689f
C2302 a_11940_14040# VSS 1.57458f
C2303 a_11654_13722# VSS 0.18412f
C2304 sg13_a21o_1_0.X VSS 1.01442f
C2305 a_11464_13854# VSS 0.10225f $ **FLOATING
C2306 a_9728_13644# VSS 0.01015f $ **FLOATING
C2307 a_11914_13945# VSS 0.24067f
C2308 a_9728_13854# VSS 0.04605f $ **FLOATING
C2309 a_8776_13644# VSS 0.02767f $ **FLOATING
C2310 a_8776_13854# VSS 0.10459f $ **FLOATING
C2311 sg13_buf_1_6.X VSS 0.70151f
C2312 a_8968_13760# VSS 0.38272f
C2313 a_25768_14570# VSS 0.12848f $ **FLOATING
C2314 a_16294_14484# VSS 0.02632f
C2315 a_25768_14914# VSS 0.02373f $ **FLOATING
C2316 a_16430_14832# VSS 0.01108f
C2317 sg13_dfrbpq_1_1.Q VSS 0.79056f
C2318 a_15784_14570# VSS 0.08916f $ **FLOATING
C2319 a_16051_14746# VSS 0.50965f
C2320 a_15784_14914# VSS 0.02464f $ **FLOATING
C2321 sg13_buf_1_0.A VSS 3.14746f
C2322 a_14098_14922# VSS 0.00329f
C2323 a_13585_14845# VSS 0.09495f
C2324 a_14346_14484# VSS 0.42699f
C2325 a_13679_14845# VSS 0.52303f
C2326 a_13936_14726# VSS 0.242f
C2327 a_12939_14495# VSS 0.36916f
C2328 a_13297_14837# VSS 0.00443f
C2329 a_12708_14909# VSS 0.03599f
C2330 a_12837_14495# VSS 0.77686f
C2331 a_12420_14488# VSS 1.57543f
C2332 a_12394_14452# VSS 0.23774f
C2333 a_12228_14922# VSS 0
C2334 a_12134_14922# VSS 0.20348f
C2335 a_17696_15156# VSS 0.00892f $ **FLOATING
C2336 a_17696_15366# VSS 0.04724f $ **FLOATING
C2337 a_16832_15156# VSS 0.00765f $ **FLOATING
C2338 sg13_a21o_1_1.A2 VSS 1.21093f
C2339 a_16832_15366# VSS 0.04127f $ **FLOATING
C2340 a_16210_15234# VSS 0.00329f
C2341 a_15697_15311# VSS 0.09495f
C2342 a_15409_15255# VSS 0.00443f
C2343 a_14820_15247# VSS 0.03599f
C2344 a_17800_15272# VSS 0.37997f
C2345 a_16458_15532# VSS 0.41936f
C2346 a_16048_15454# VSS 0.2428f
C2347 a_15791_15311# VSS 0.5218f
C2348 a_14340_15234# VSS 0
C2349 a_11848_15156# VSS 0.02614f $ **FLOATING
C2350 a_15051_15356# VSS 0.37179f
C2351 a_14949_15213# VSS 0.78001f
C2352 a_14532_15552# VSS 1.57404f
C2353 a_14246_15234# VSS 0.17239f
C2354 sg13_dfrbpq_1_3.D VSS 0.61189f
C2355 a_14506_15457# VSS 0.23687f
C2356 a_12650_15532# VSS 0
C2357 sg13_nor2b_1_0.Y VSS 0.54646f
C2358 a_12268_15532# VSS 0
C2359 a_11848_15366# VSS 0.08318f $ **FLOATING
C2360 a_12046_15276# VSS 0.36098f
C2361 a_16735_15972# VSS 0.00152f
C2362 a_17006_16388# VSS 0.00578f
C2363 sg13_inv_1_1.A VSS 0.42413f
C2364 a_16018_16434# VSS 0.00329f
C2365 a_15505_16357# VSS 0.09498f
C2366 sg13_inv_2_1.A VSS 1.40789f
C2367 sg13_dfrbpq_1_3.Q VSS 1.2999f
C2368 a_16266_15996# VSS 0.41808f
C2369 a_15599_16357# VSS 0.52252f
C2370 a_15856_16238# VSS 0.24086f
C2371 a_14859_16007# VSS 0.37055f
C2372 a_15217_16349# VSS 0.00443f
C2373 a_14628_16421# VSS 0.03599f
C2374 a_13864_16082# VSS 0.08174f $ **FLOATING
C2375 a_13499_15996# VSS 0.00632f
C2376 a_14757_16007# VSS 0.78589f
C2377 a_14340_16000# VSS 1.57504f
C2378 a_14314_15964# VSS 0.2373f
C2379 a_14148_16434# VSS 0
C2380 a_14054_16434# VSS 0.18236f
C2381 sg13_inv_1_1.Y VSS 0.342f
C2382 a_13864_16426# VSS 0.0234f $ **FLOATING
C2383 a_13601_16344# VSS 0.01118f
C2384 sg13_nor2_1_0.Y VSS 0.66093f
C2385 sg13_nor2_1_0.B VSS 0.93284f
C2386 a_12754_16434# VSS 0.00329f
C2387 a_12241_16357# VSS 0.09499f
C2388 a_13002_15996# VSS 0.42042f
C2389 a_12335_16357# VSS 0.52459f
C2390 a_12592_16238# VSS 0.23909f
C2391 a_11595_16007# VSS 0.37009f
C2392 a_11953_16349# VSS 0.00443f
C2393 a_11364_16421# VSS 0.03599f
C2394 a_11493_16007# VSS 0.77341f
C2395 a_11076_16000# VSS 1.57798f
C2396 a_11050_15964# VSS 0.23857f
C2397 a_10884_16434# VSS 0
C2398 a_10790_16434# VSS 0.20578f
C2399 sg13_dfrbpq_1_4.D VSS 0.3693f
C2400 sg13_nor2_1_0.A VSS 1.02565f
C2401 a_9920_16082# VSS 0.04735f $ **FLOATING
C2402 a_10024_15996# VSS 0.37713f
C2403 a_9920_16426# VSS 0.00892f $ **FLOATING
C2404 a_7816_15996# VSS 0.38385f
C2405 a_25856_16668# VSS 0.00748f $ **FLOATING
C2406 a_25856_16878# VSS 0.08592f $ **FLOATING
C2407 a_15680_16668# VSS 0.00697f $ **FLOATING
C2408 a_15496_16668# VSS 0.01913f $ **FLOATING
C2409 a_15680_16878# VSS 0.03558f $ **FLOATING
C2410 a_15496_16878# VSS 0.0819f $ **FLOATING
C2411 a_14912_16668# VSS 0.0054f $ **FLOATING
C2412 a_14998_16742# VSS 0.22026f
C2413 sg13_dfrbpq_1_5.Q VSS 1.1949f
C2414 a_14912_16878# VSS 0.0424f $ **FLOATING
C2415 a_14290_16746# VSS 0.00329f
C2416 a_13777_16823# VSS 0.095f
C2417 a_13489_16767# VSS 0.00443f
C2418 a_12900_16759# VSS 0.03599f
C2419 sg13_o21ai_1_0.A1 VSS 0.5681f
C2420 a_14538_17044# VSS 0.41947f
C2421 a_14128_16966# VSS 0.2437f
C2422 a_13871_16823# VSS 0.51719f
C2423 a_12420_16746# VSS 0
C2424 a_12136_16668# VSS 0.02444f $ **FLOATING
C2425 sg13_dfrbpq_1_0.CLK VSS 3.32437f
C2426 a_13131_16868# VSS 0.37453f
C2427 a_13029_16725# VSS 0.79298f
C2428 a_12612_17064# VSS 1.57631f
C2429 a_12326_16746# VSS 0.18395f
C2430 sg13_dfrbpq_1_6.D VSS 0.5976f
C2431 a_12136_16878# VSS 0.1023f $ **FLOATING
C2432 sg13_inv_1_0.Y VSS 6.6032f
C2433 a_12586_16969# VSS 0.24067f
C2434 a_25856_17594# VSS 0.08592f $ **FLOATING
C2435 a_25856_17938# VSS 0.00748f $ **FLOATING
C2436 sg13_o21ai_1_0.B1 VSS 0.57643f
C2437 a_14437_17878# VSS 0.00852f
C2438 a_14144_17594# VSS 0.05786f $ **FLOATING
C2439 a_14235_17564# VSS 0.38895f
C2440 a_14144_17938# VSS 0.00899f $ **FLOATING
C2441 a_25768_23642# VSS 0.12888f $ **FLOATING
C2442 a_25768_23986# VSS 0.02422f $ **FLOATING
C2443 a_14144_23642# VSS 0.06023f $ **FLOATING
C2444 sg13_a21oi_1_0.A1 VSS 2.2072f
C2445 a_14248_23556# VSS 0.38693f
C2446 a_14144_23986# VSS 0.00902f $ **FLOATING
C2447 a_25768_25154# VSS 0.14597f $ **FLOATING
C2448 a_25768_25498# VSS 0.02451f $ **FLOATING
C2449 sg13_a22oi_1_0.B2 VSS 3.0457f
C2450 a_15872_25154# VSS 0.03985f $ **FLOATING
C2451 a_15688_25154# VSS 0.10206f $ **FLOATING
C2452 a_15976_25068# VSS 0.384f
C2453 a_15872_25498# VSS 0.00693f $ **FLOATING
C2454 a_15688_25498# VSS 0.02637f $ **FLOATING
C2455 sg13_a21oi_1_0.A2 VSS 2.71f
C2456 a_13856_25154# VSS 0.04901f $ **FLOATING
C2457 a_13960_25068# VSS 0.38011f
C2458 a_13856_25498# VSS 0.00907f $ **FLOATING
.ends

